CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 429
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 429
8912914 0
0
6 Title:
5 Name:
0
0
0
9
7 Ground~
168 128 217 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
11 Signal Gen~
195 93 179 0 24 64
0 7 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846079 0 1084227584
0 897988541 897988541 973279855 981668463
20
0 1000 0 5 0 1e-006 1e-006 0.0005 0.001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 336 0
4 0/5V
-15 -30 13 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 PULSE(0 5 0 1u 1u 500u 1m)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
4 7445
219 352 138 0 14 29
0 11 10 9 8 12 13 14 6 15
16 5 17 18 19
0
0 0 12528 0
4 7445
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 1
2 3 4 5 6 7 9 10 11 0
65 0 0 512 1 0 0 0
1 U
3618 0 0
0
0
7 74LS293
154 235 165 0 8 17
0 2 2 7 8 11 10 9 8
0
0 0 12528 0
7 74LS293
-24 -35 25 -27
2 U2
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
7 Ground~
168 174 217 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
2 +V
167 448 54 0 1 3
0 3
0
0 0 53616 0
4 +24V
-14 -15 14 -7
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7734 0 0
0
0
2 +V
167 508 76 0 1 3
0 4
0
0 0 53616 0
4 +24V
-14 -15 14 -7
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
9 Resistor~
219 448 96 0 3 5
0 3 5 1
0
0 0 112 270
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 508 120 0 3 5
0 4 6 1
0
0 0 112 270
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
13
1 1 3 0 0 4224 0 8 6 0 0 2
448 78
448 63
1 2 2 0 0 4096 0 1 2 0 0 3
128 211
128 184
124 184
1 1 4 0 0 4224 0 9 7 0 0 2
508 102
508 85
2 11 5 0 0 8320 0 8 3 0 0 3
448 114
448 129
390 129
2 8 6 0 0 8320 0 9 3 0 0 3
508 138
508 156
390 156
2 0 2 0 0 4096 0 4 0 0 7 2
203 165
174 165
1 1 2 0 0 8320 0 4 5 0 0 3
203 156
174 156
174 211
1 3 7 0 0 4224 0 2 4 0 0 2
124 174
197 174
0 4 8 0 0 8320 0 0 4 10 0 5
278 183
278 205
188 205
188 183
197 183
8 4 8 0 0 0 0 4 3 0 0 2
267 183
320 183
7 3 9 0 0 4224 0 4 3 0 0 2
267 174
320 174
6 2 10 0 0 4224 0 4 3 0 0 2
267 165
320 165
5 1 11 0 0 4224 0 4 3 0 0 2
267 156
320 156
1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 80
110 254 470 298
114 258 466 290
80 Counter/decoder combination used to provide 
timing and sequencing operations.
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.016 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
296681548 8525888 100 100 0 0
77 66 587 216
4 430 635 712
530 66
77 66
587 141
587 141
0 0
0.0159882 0 0 0 0.016 0.016
13425 0
2 0.003 20
3
150 174
0 7 0 50 1	0 8 0 0
419 156
0 6 0 0 2	0 5 0 0
421 129
0 5 0 -50 2	0 4 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
9.98039 0 5.4 0 10 10
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 14 0 0
200 112
0 7 0 0 2	0 14 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
