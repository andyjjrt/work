CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 432
8388626 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 150 54 0 1 11
0 5
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
1 A
-24 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 150 89 0 1 11
0 4
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
1 B
-23 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 150 131 0 1 11
0 3
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
3 Cin
-37 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
14 Logic Display~
6 442 50 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
5 4081~
219 289 145 0 3 22
0 4 3 8
0
0 0 96 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
5394 0 0
0
0
5 4081~
219 289 192 0 3 22
0 4 5 7
0
0 0 96 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
7734 0 0
0
0
5 4081~
219 289 238 0 3 22
0 3 5 6
0
0 0 96 0
4 4081
-7 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 1 0
1 U
9914 0 0
0
0
5 4030~
219 360 76 0 3 22
0 5 10 11
0
0 0 96 0
4 4030
-7 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 2 0
1 U
3747 0 0
0
0
5 4030~
219 281 98 0 3 22
0 4 3 10
0
0 0 96 0
4 4030
-7 -24 21 -16
3 U2B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
3549 0 0
0
0
8 3-In OR~
219 360 192 0 4 22
0 8 7 6 9
0
0 0 96 0
4 4075
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 3 0
1 U
7931 0 0
0
0
14 Logic Display~
6 442 161 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
16
0 0 2 0 0 12672 0 0 0 0 0 6
180 31
180 275
410 275
410 27
180 27
180 31
0 1 3 0 0 4096 0 0 3 8 0 2
229 131
162 131
1 0 4 0 0 4096 0 5 0 0 7 2
265 136
247 136
2 0 3 0 0 0 0 5 0 0 8 2
265 154
229 154
2 0 5 0 0 4096 0 6 0 0 6 2
265 201
213 201
2 0 5 0 0 8320 0 7 0 0 15 3
265 247
213 247
213 54
1 0 4 0 0 8192 0 6 0 0 9 3
265 183
247 183
247 89
1 2 3 0 0 8320 0 7 9 0 0 4
265 229
229 229
229 107
265 107
1 1 4 0 0 4224 0 9 2 0 0 2
265 89
162 89
3 3 6 0 0 8320 0 10 7 0 0 4
347 201
335 201
335 238
310 238
2 3 7 0 0 4224 0 10 6 0 0 2
348 192
310 192
1 3 8 0 0 8320 0 10 5 0 0 4
347 183
335 183
335 145
310 145
4 1 9 0 0 4224 0 10 11 0 0 3
393 192
442 192
442 179
2 3 10 0 0 12416 0 8 9 0 0 4
344 85
335 85
335 98
314 98
1 1 5 0 0 0 0 8 1 0 0 4
344 67
335 67
335 54
162 54
1 3 11 0 0 8320 0 4 8 0 0 3
442 68
442 76
393 76
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 36
150 288 446 312
154 292 442 308
36 Complete circuitry for a full adder.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
422 190 462 214
426 194 458 210
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
435 74 451 98
439 78 447 94
1 S
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
