CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 534
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 534
8388626 0
0
6 Title:
5 Name:
0
0
0
44
14 Logic Display~
6 175 36 0 1 2
10 2
0
0 0 54384 0
6 100MEG
3 -16 45 -8
3 L24
-11 -21 10 -13
1 A
-4 -21 3 -13
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8953 0 0
0
0
14 Logic Display~
6 164 36 0 1 2
10 3
0
0 0 54384 0
6 100MEG
3 -16 45 -8
3 L23
-11 -21 10 -13
1 B
-4 -21 3 -13
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 153 36 0 1 2
10 4
0
0 0 54384 0
6 100MEG
3 -16 45 -8
3 L22
-11 -21 10 -13
1 C
-4 -21 3 -13
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 142 36 0 1 2
10 5
0
0 0 54384 0
6 100MEG
3 -16 45 -8
3 L21
-11 -21 10 -13
1 D
-4 -21 3 -13
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
6 74LS42
101 514 148 0 14 29
0 5 4 3 2 10 12 11 13 14
15 16 17 18 19
0
0 0 5232 270
6 74LS42
-21 -60 21 -52
2 U8
60 -5 74 3
4 7442
-11 -5 17 3
15 DVCC=16;DGND=8;
106 %D [%16bi %8bi %1i %2i %3i %4i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 11 10 9 7 6
5 4 3 2 1 12 13 14 15 11
10 9 7 6 5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
5394 0 0
0
0
14 Logic Display~
6 330 304 0 1 2
10 37
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
9 Inverter~
13 351 136 0 2 22
0 5 35
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U6B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 6 0
1 U
9914 0 0
0
0
9 Inverter~
13 351 180 0 2 22
0 35 36
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U6A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
3747 0 0
0
0
10 4-In NAND~
219 61 265 0 5 22
0 20 33 34 35 23
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U1A
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 1 0
1 U
3549 0 0
0
0
10 4-In NAND~
219 100 265 0 5 22
0 33 34 35 32 24
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U1B
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 1 0
1 U
7931 0 0
0
0
10 4-In NAND~
219 138 265 0 5 22
0 35 34 20 21 27
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U2A
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 2 0
1 U
9325 0 0
0
0
10 4-In NAND~
219 176 265 0 5 22
0 35 21 34 32 26
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U2B
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 2 0
1 U
8903 0 0
0
0
10 4-In NAND~
219 214 265 0 5 22
0 35 33 22 20 25
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U3A
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 3 0
1 U
3834 0 0
0
0
10 4-In NAND~
219 405 265 0 5 22
0 32 33 34 36 30
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U3B
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 3 0
1 U
3363 0 0
0
0
10 4-In NAND~
219 367 265 0 5 22
0 20 33 34 36 31
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U4A
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
7668 0 0
0
0
10 4-In NAND~
219 329 265 0 5 22
0 32 21 22 35 37
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U4B
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 4 0
1 U
4718 0 0
0
0
10 4-In NAND~
219 291 265 0 5 22
0 35 20 21 22 29
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U5A
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 5 0
1 U
3874 0 0
0
0
10 4-In NAND~
219 252 265 0 5 22
0 35 33 32 22 28
0
0 0 112 270
6 74LS20
-21 -28 21 -20
3 U5B
22 -7 43 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 5 0
1 U
6671 0 0
0
0
9 Inverter~
13 269 179 0 2 22
0 34 22
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U6C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 6 0
1 U
3789 0 0
0
0
9 Inverter~
13 269 136 0 2 22
0 4 34
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U6D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 6 0
1 U
4871 0 0
0
0
9 Inverter~
13 193 179 0 2 22
0 33 21
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U6E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 6 0
1 U
3750 0 0
0
0
9 Inverter~
13 193 136 0 2 22
0 3 33
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U6F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 6 0
1 U
8778 0 0
0
0
9 Inverter~
13 116 179 0 2 22
0 20 32
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U7A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
538 0 0
0
0
9 Inverter~
13 116 136 0 2 22
0 2 20
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U7B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 7 0
1 U
6843 0 0
0
0
14 Logic Display~
6 368 304 0 1 2
10 31
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3136 0 0
0
0
14 Logic Display~
6 406 304 0 1 2
10 30
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5950 0 0
0
0
14 Logic Display~
6 292 304 0 1 2
10 29
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
14 Logic Display~
6 253 304 0 1 2
10 28
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6828 0 0
0
0
14 Logic Display~
6 62 304 0 1 2
10 23
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
14 Logic Display~
6 101 304 0 1 2
10 24
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L7
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8365 0 0
0
0
14 Logic Display~
6 215 304 0 1 2
10 25
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L8
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4132 0 0
0
0
14 Logic Display~
6 177 304 0 1 2
10 26
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4551 0 0
0
0
14 Logic Display~
6 139 304 0 1 2
10 27
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L10
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3635 0 0
0
0
9 Data Seq~
170 73 55 0 17 18
0 39 40 41 42 5 4 3 2 43
44 15 1 16 5 1 0 33
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
3973 0 0
0
0
AAAAABACADAEAFAGAHAIAJAKALAMANAOAPAAABACADAEAFAGAHAIAJAKALAMANAOAP
14 Logic Display~
6 474 198 0 1 2
10 19
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L11
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3851 0 0
0
0
14 Logic Display~
6 483 198 0 1 2
10 18
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L12
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8383 0 0
0
0
14 Logic Display~
6 501 198 0 1 2
10 16
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L13
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9334 0 0
0
0
14 Logic Display~
6 492 198 0 1 2
10 17
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L14
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7471 0 0
0
0
14 Logic Display~
6 510 198 0 1 2
10 15
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L15
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3334 0 0
0
0
14 Logic Display~
6 555 198 0 1 2
10 10
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L16
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3559 0 0
0
0
14 Logic Display~
6 537 198 0 1 2
10 11
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L17
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
984 0 0
0
0
14 Logic Display~
6 546 198 0 1 2
10 12
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L18
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7557 0 0
0
0
14 Logic Display~
6 528 198 0 1 2
10 13
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L19
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3146 0 0
0
0
14 Logic Display~
6 519 198 0 1 2
10 14
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L20
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5687 0 0
0
0
80
1 0 2 0 0 4096 0 1 0 0 12 2
175 54
175 91
1 0 3 0 0 4096 0 2 0 0 28 2
164 54
164 82
1 0 4 0 0 4096 0 3 0 0 27 2
153 54
153 73
1 0 5 0 0 4096 0 4 0 0 26 2
142 54
142 64
0 0 6 0 0 4224 0 0 0 0 0 2
441 150
456 150
0 0 7 0 0 4224 0 0 0 0 0 2
441 146
456 146
0 0 8 0 0 4224 0 0 0 0 0 2
441 142
456 142
0 0 9 0 0 4480 0 0 0 0 0 5
37 285
430 285
430 112
37 112
37 276
0 1 5 0 0 4096 0 0 5 26 0 3
354 64
501 64
501 115
0 2 4 0 0 4224 0 0 5 27 0 3
272 73
492 73
492 115
0 3 3 0 0 4224 0 0 5 28 0 3
196 82
483 82
483 115
0 4 2 0 0 4224 0 0 5 29 0 3
119 91
474 91
474 115
1 5 10 0 0 4224 0 40 5 0 0 2
555 184
555 185
1 7 11 0 0 4224 0 41 5 0 0 2
537 184
537 185
1 6 12 0 0 4224 0 42 5 0 0 2
546 184
546 185
1 8 13 0 0 4224 0 43 5 0 0 2
528 184
528 185
1 9 14 0 0 4224 0 44 5 0 0 2
519 184
519 185
1 10 15 0 0 4224 0 39 5 0 0 2
510 184
510 185
1 11 16 0 0 4224 0 37 5 0 0 2
501 184
501 185
1 12 17 0 0 4224 0 38 5 0 0 2
492 184
492 185
1 13 18 0 0 4224 0 36 5 0 0 2
483 184
483 185
1 14 19 0 0 4224 0 35 5 0 0 2
474 184
474 185
2 0 20 0 0 4096 0 17 0 0 72 2
296 240
296 207
3 0 21 0 0 4096 0 17 0 0 73 2
287 240
287 212
4 0 22 0 0 4096 0 17 0 0 75 2
278 240
278 222
5 1 5 0 0 4224 0 34 7 0 0 3
105 64
354 64
354 118
6 1 4 0 0 0 0 34 20 0 0 3
105 73
272 73
272 118
7 1 3 0 0 0 0 34 22 0 0 3
105 82
196 82
196 118
8 1 2 0 0 0 0 34 24 0 0 3
105 91
119 91
119 118
1 5 23 0 0 4224 0 29 9 0 0 2
62 290
62 291
1 5 24 0 0 4224 0 30 10 0 0 2
101 290
101 291
1 5 25 0 0 4224 0 31 13 0 0 2
215 290
215 291
1 5 26 0 0 4224 0 32 12 0 0 2
177 290
177 291
1 5 27 0 0 4224 0 33 11 0 0 2
139 290
139 291
1 5 28 0 0 4224 0 28 18 0 0 2
253 290
253 291
1 5 29 0 0 4224 0 27 17 0 0 2
292 290
292 291
1 5 30 0 0 4224 0 26 14 0 0 2
406 290
406 291
1 5 31 0 0 4224 0 25 15 0 0 2
368 290
368 291
0 0 20 0 0 4096 0 0 0 72 62 3
75 207
75 157
119 157
2 0 32 0 0 4096 0 23 0 0 71 2
119 197
119 202
1 0 33 0 0 4096 0 10 0 0 74 2
114 240
114 217
2 0 34 0 0 4096 0 10 0 0 76 2
105 240
105 227
3 0 35 0 0 4096 0 10 0 0 77 2
96 240
96 232
0 0 33 0 0 4096 0 0 0 74 63 3
158 217
158 158
196 158
3 0 20 0 0 0 0 11 0 0 72 2
134 240
134 207
2 0 34 0 0 0 0 11 0 0 76 2
143 240
143 227
1 0 35 0 0 0 0 11 0 0 77 2
152 240
152 232
4 0 32 0 0 4096 0 12 0 0 71 2
163 240
163 202
3 0 34 0 0 0 0 12 0 0 76 2
172 240
172 227
2 0 21 0 0 0 0 12 0 0 73 2
181 240
181 212
1 0 35 0 0 0 0 12 0 0 77 2
190 240
190 232
2 0 21 0 0 0 0 21 0 0 73 2
196 197
196 212
4 0 20 0 0 0 0 13 0 0 72 2
201 240
201 207
0 0 34 0 0 8192 0 0 0 64 76 3
272 157
233 157
233 227
2 0 33 0 0 0 0 13 0 0 74 2
219 240
219 217
1 0 35 0 0 0 0 13 0 0 77 2
228 240
228 232
4 0 22 0 0 0 0 18 0 0 75 2
239 240
239 222
3 0 32 0 0 0 0 18 0 0 71 2
248 240
248 202
2 0 33 0 0 0 0 18 0 0 74 2
257 240
257 217
1 0 35 0 0 0 0 18 0 0 77 2
266 240
266 232
2 0 22 0 0 4096 0 19 0 0 75 2
272 197
272 222
2 1 20 0 0 0 0 24 23 0 0 2
119 154
119 161
2 1 33 0 0 0 0 22 21 0 0 2
196 154
196 161
2 1 34 0 0 0 0 20 19 0 0 2
272 154
272 161
1 0 35 0 0 0 0 17 0 0 77 2
305 240
305 232
1 0 32 0 0 0 0 16 0 0 71 2
343 240
343 202
2 1 35 0 0 0 0 7 8 0 0 2
354 154
354 162
0 0 35 0 0 4096 0 0 0 77 67 3
316 232
316 157
354 157
2 0 33 0 0 0 0 15 0 0 74 2
372 240
372 217
3 0 34 0 0 0 0 15 0 0 76 2
363 240
363 227
1 4 32 0 0 8320 0 14 10 0 0 4
419 240
419 202
87 202
87 240
1 1 20 0 0 8320 0 15 9 0 0 4
381 240
381 207
75 207
75 240
2 4 21 0 0 8320 0 16 11 0 0 4
334 240
334 212
125 212
125 240
2 2 33 0 0 8320 0 14 9 0 0 4
410 240
410 217
66 217
66 240
3 3 22 0 0 8320 0 16 13 0 0 4
325 240
325 222
210 222
210 240
3 3 34 0 0 8320 0 14 9 0 0 4
401 240
401 227
57 227
57 240
4 4 35 0 0 8320 0 16 9 0 0 4
316 240
316 232
48 232
48 240
4 0 36 0 0 8192 0 14 0 0 79 3
392 240
392 232
354 232
2 4 36 0 0 4224 0 8 15 0 0 2
354 198
354 240
1 5 37 0 0 4224 0 6 16 0 0 2
330 290
330 291
29
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 50
104 386 512 410
108 390 508 406
50 Logic diagram for the 7442 BCD-to-decimal decoder.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
36 110 71 130
40 114 68 128
4 7442
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
50 319 71 339
54 323 68 337
2 O0
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
50 307 64 327
54 311 61 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
90 307 104 327
94 311 101 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
90 319 111 339
94 323 108 337
2 O1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
129 319 150 339
133 323 147 337
2 O2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
166 319 187 339
170 323 184 337
2 O3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
204 319 225 339
208 323 222 337
2 O4
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
242 319 263 339
246 323 260 337
2 O5
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
281 319 302 339
285 323 299 337
2 O6
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
319 319 340 339
323 323 337 337
2 O7
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
357 319 378 339
361 323 375 337
2 O8
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
396 319 417 339
400 323 414 337
2 O9
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
129 307 143 327
133 311 140 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
166 307 180 327
170 311 177 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
204 307 218 327
208 311 215 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
242 307 256 327
246 311 253 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
281 307 295 327
285 311 292 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
319 307 333 327
323 311 330 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
357 307 371 327
361 311 368 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
396 307 410 327
400 311 407 325
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
462 212 567 232
466 216 564 230
14 O0----------O9
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
462 200 476 220
466 204 473 218
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
546 200 560 220
550 204 557 218
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
119 94 133 114
123 98 130 112
1 A
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
196 94 210 114
200 98 207 112
1 B
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
271 94 285 114
275 98 282 112
1 C
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
353 93 367 113
357 97 364 111
1 D
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
267780172 8525888 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
9.98039 0 5.4 0 10 10
12401 0
4 1e-006 2
2
221 112
0 7 0 0 2	0 81 0 0
367 106
0 2 0 0 1	0 81 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 81 0 0
200 112
0 7 0 0 2	0 81 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
