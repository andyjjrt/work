CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 395
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 395 635 522
25165842 0
0
6 Title:
5 Name:
0
0
0
8
7 Ground~
168 229 74 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
7 Ground~
168 243 157 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
5 SCOPE
12 128 90 0 1 11
0 6
0
0 0 57568 0
1 J
-4 -4 3 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 163 90 0 1 11
0 5
0
0 0 57568 0
1 K
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
5 SCOPE
12 198 90 0 1 11
0 4
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 286 91 0 1 11
0 7
0
0 0 57568 0
1 Q
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
9 Data Seq~
170 72 92 0 17 18
0 11 12 13 14 15 6 4 5 16
17 6 5 50 2 1 0 51
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
9914 0 0
0
0
AAAAAAACACAAABADAHAFAFAHACAAAAACAGAEAEAGAHAFAFAHAHAFAFAHIHAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAA
5 4027~
219 243 146 0 7 32
0 2 6 4 5 2 18 7
0
0 0 4192 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 512 2 1 6 0
1 U
3747 0 0
0
0
14
0 0 3 0 0 16 0 0 0 0 0 5
320 232
592 232
592 264
320 264
320 232
1 1 2 0 0 12416 0 1 8 0 0 4
229 68
229 64
243 64
243 89
1 5 2 0 0 0 0 2 8 0 0 2
243 151
243 152
1 0 4 0 0 4096 0 5 0 0 9 2
198 102
198 119
1 0 5 0 0 4096 0 4 0 0 8 2
163 102
163 128
1 0 6 0 0 4096 0 3 0 0 10 2
128 102
128 110
1 7 7 0 0 8320 0 6 8 0 0 3
286 103
286 110
267 110
8 4 5 0 0 4224 0 7 8 0 0 2
104 128
219 128
7 3 4 0 0 4224 0 7 8 0 0 2
104 119
219 119
6 2 6 0 0 4224 0 7 8 0 0 2
104 110
219 110
0 0 1 0 0 4256 0 0 0 12 14 2
436 64
436 148
0 0 8 0 0 4224 0 0 0 0 0 2
342 64
563 64
0 0 9 0 0 4224 0 0 0 0 0 2
342 80
563 80
0 0 10 0 0 4224 0 0 0 0 0 2
342 148
563 148
15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 81
24 217 280 281
28 221 276 269
81 Clocked J-K flip-flop that 
responds only to the positive 
edge of the clock.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
322 229 588 266
326 233 585 261
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 43
441 61 569 165
445 65 565 145
43       Q
Qo (no change)
1
0
Qo (toggles)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
403 95 419 119
407 99 415 115
1 ^
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
403 93 419 117
407 97 415 113
1 |
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
396 61 428 85
400 65 424 81
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
403 125 419 149
407 129 415 145
1 |
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
403 127 419 151
407 131 415 147
1 ^
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
403 110 419 134
407 114 415 130
1 |
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
403 112 419 136
407 116 415 132
1 ^
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
403 75 419 99
407 79 415 95
1 |
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
403 77 419 101
407 81 415 97
1 ^
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
349 61 373 165
353 65 369 145
13 J
0
1
0
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
376 61 400 165
380 65 396 145
13 K
0
0
1
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
441 111 465 135
445 115 461 131
2 __
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 4.6e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
