CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 435
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 435 635 561
25165842 0
0
6 Title:
5 Name:
0
0
0
33
13 Logic Switch~
5 409 260 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21600 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
7 Up/Down
-66 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
9 Inverter~
13 485 217 0 2 22
0 14 13
0
0 0 96 512
6 74LS04
-21 -19 21 -11
3 U6A
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 6 0
1 U
4441 0 0
0
0
5 4081~
219 421 123 0 3 22
0 14 2 19
0
0 0 1120 512
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
1 1
-4 -5 3 3
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
3618 0 0
0
0
5 4073~
219 232 107 0 4 22
0 14 2 4 16
0
0 0 1120 512
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
1 2
-4 -5 3 3
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 2 0
1 U
6153 0 0
0
0
5 4081~
219 423 191 0 3 22
0 3 13 20
0
0 0 1120 512
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
1 3
-4 -5 3 3
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
5394 0 0
0
0
5 4073~
219 232 208 0 4 22
0 18 3 13 17
0
0 0 1120 512
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
1 4
-4 -5 3 3
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 2 0
1 U
7734 0 0
0
0
5 4071~
219 369 157 0 3 22
0 19 20 15
0
0 0 96 512
4 4071
-7 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 5 0
1 U
9914 0 0
0
0
5 4071~
219 171 157 0 3 22
0 16 17 12
0
0 0 96 512
4 4071
-7 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 5 0
1 U
3747 0 0
0
0
6 74113~
219 485 165 0 6 22
0 11 8 11 11 3 2
0
0 0 4192 512
7 74LS113
-25 -42 24 -34
3 U4A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 1 4 0
1 U
3549 0 0
0
0
6 74113~
219 296 165 0 6 22
0 15 8 15 10 18 4
0
0 0 4192 512
7 74LS113
-25 -42 24 -34
3 U4B
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 2 4 0
1 U
7931 0 0
0
0
6 74113~
219 100 165 0 6 22
0 12 8 12 9 21 5
0
0 0 4192 512
7 74LS113
-25 -42 24 -34
3 U3A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 3 0
1 U
9325 0 0
0
0
7 Pulser~
4 80 223 0 10 12
0 22 23 8 24 0 0 5 5 6
7
0
0 0 5152 0
0
2 V2
-7 -28 7 -20
5 CLOCK
-18 -28 17 -20
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8903 0 0
0
0
2 +V
167 483 116 0 1 3
0 11
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
0
0
9 Terminal~
194 269 108 0 1 3
0 2
0
0 0 49504 270
1 A
2 -5 9 3
2 T3
-7 -32 7 -24
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3363 0 0
0
0
9 Terminal~
194 438 150 0 1 3
0 2
0
0 0 49504 90
1 A
-10 -5 -3 3
2 T1
-7 -32 7 -24
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7668 0 0
0
0
9 Terminal~
194 439 168 0 1 3
0 3
0
0 0 49504 90
2 AN
-19 -5 -5 3
2 T2
-7 -32 7 -24
0
3 AN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4718 0 0
0
0
9 Terminal~
194 271 209 0 1 3
0 3
0
0 0 49504 270
2 AN
2 -5 16 3
2 T4
-7 -32 7 -24
0
3 AN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3874 0 0
0
0
2 +V
167 294 114 0 1 3
0 10
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6671 0 0
0
0
2 +V
167 98 115 0 1 3
0 9
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3789 0 0
0
0
9 Terminal~
194 243 150 0 1 3
0 4
0
0 0 49504 90
1 B
-9 -6 -2 2
2 T5
-7 -25 7 -17
0
2 B;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4871 0 0
0
0
9 Terminal~
194 60 150 0 1 3
0 5
0
0 0 49504 90
1 C
-11 -6 -4 2
2 T6
-7 -25 7 -17
0
2 C;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3750 0 0
0
0
5 SCOPE
12 166 229 0 1 11
0 8
0
0 0 57568 0
2 CP
-8 -4 6 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8778 0 0
0
0
9 Terminal~
194 163 78 0 1 3
0 2
0
0 0 49504 180
1 A
6 -7 13 1
2 T9
3 -17 17 -9
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
538 0 0
0
0
9 Terminal~
194 112 83 0 1 3
0 4
0
0 0 49504 180
1 B
6 -7 13 1
2 T8
3 -17 17 -9
0
2 B;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6843 0 0
0
0
9 Terminal~
194 61 88 0 1 3
0 5
0
0 0 49504 180
1 C
6 -7 13 1
2 T7
3 -17 17 -9
0
2 C;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3136 0 0
0
0
7 Ground~
168 15 103 0 1 3
0 6
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5950 0 0
0
0
14 Logic Display~
6 186 19 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
5 SCOPE
12 163 25 0 1 11
0 2
0
0 0 57568 0
1 A
-4 -4 3 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6828 0 0
0
0
14 Logic Display~
6 135 19 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
5 SCOPE
12 112 25 0 1 11
0 4
0
0 0 57568 0
1 B
-4 -4 3 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8365 0 0
0
0
14 Logic Display~
6 84 19 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4132 0 0
0
0
5 SCOPE
12 61 25 0 1 11
0 5
0
0 0 57568 0
1 C
-4 -4 3 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4551 0 0
0
0
12 Hex Display~
7 24 35 0 16 19
10 2 4 5 6 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3635 0 0
0
0
43
0 0 7 0 0 4240 0 0 0 0 0 5
304 11
575 11
575 44
304 44
304 11
1 0 8 0 0 0 0 22 0 0 28 2
166 241
166 241
1 6 5 0 0 4096 0 21 11 0 0 2
71 148
74 148
1 0 4 0 0 0 0 20 0 0 17 2
254 148
254 148
1 4 9 0 0 4224 0 19 11 0 0 2
98 124
98 121
1 4 10 0 0 4224 0 18 10 0 0 2
294 123
294 121
1 2 3 0 0 4096 0 17 6 0 0 2
259 208
252 208
1 2 2 0 0 4096 0 14 4 0 0 2
257 107
252 107
1 0 3 0 0 0 0 16 0 0 32 2
450 166
449 166
1 0 2 0 0 0 0 15 0 0 33 2
449 148
449 148
1 0 11 0 0 4096 0 9 0 0 12 2
507 148
526 148
0 3 11 0 0 4224 0 0 9 13 0 4
483 123
526 123
526 166
507 166
1 4 11 0 0 0 0 13 9 0 0 2
483 125
483 121
3 0 8 0 0 8192 0 12 0 0 28 4
104 214
117 214
117 241
128 241
3 0 12 0 0 4096 0 8 0 0 16 2
144 157
138 157
1 3 12 0 0 8320 0 11 11 0 0 4
122 148
138 148
138 166
122 166
6 3 4 0 0 8192 0 10 4 0 0 4
270 148
254 148
254 116
252 116
2 0 13 0 0 8192 0 5 0 0 25 3
443 200
449 200
449 217
1 0 14 0 0 8192 0 3 0 0 26 3
441 114
449 114
449 98
3 0 15 0 0 4096 0 7 0 0 29 2
342 157
335 157
4 1 16 0 0 8320 0 4 8 0 0 4
207 107
201 107
201 148
190 148
4 2 17 0 0 8320 0 6 8 0 0 4
207 208
201 208
201 166
190 166
5 1 18 0 0 8320 0 10 6 0 0 4
264 166
254 166
254 199
252 199
1 0 14 0 0 4096 0 2 0 0 26 2
506 217
540 217
3 2 13 0 0 4224 0 6 2 0 0 2
252 217
470 217
1 1 14 0 0 4224 0 4 1 0 0 4
252 98
540 98
540 260
421 260
2 0 8 0 0 4096 0 10 0 0 28 2
325 157
325 241
2 2 8 0 0 12416 0 9 11 0 0 6
514 157
517 157
517 241
128 241
128 157
129 157
1 3 15 0 0 8320 0 10 10 0 0 4
318 148
335 148
335 166
318 166
3 1 19 0 0 4224 0 3 7 0 0 3
396 123
396 148
388 148
3 2 20 0 0 8320 0 5 7 0 0 4
398 191
396 191
396 166
388 166
5 1 3 0 0 8320 0 9 5 0 0 4
453 166
449 166
449 182
443 182
6 2 2 0 0 8192 0 9 3 0 0 4
459 148
449 148
449 132
441 132
1 0 2 0 0 0 0 23 0 0 43 2
163 63
163 63
1 0 4 0 0 0 0 24 0 0 42 2
112 68
112 68
1 0 5 0 0 0 0 25 0 0 41 2
61 73
61 73
1 4 6 0 0 4224 0 26 33 0 0 2
15 97
15 59
1 0 5 0 0 4096 0 31 0 0 41 2
84 37
61 37
1 0 4 0 0 0 0 29 0 0 42 2
135 37
112 37
1 0 2 0 0 4096 0 27 0 0 43 2
186 37
163 37
3 1 5 0 0 8320 0 33 32 0 0 4
21 59
21 73
61 73
61 37
2 1 4 0 0 8320 0 33 30 0 0 4
27 59
27 68
112 68
112 37
1 1 2 0 0 8320 0 33 28 0 0 4
33 59
33 63
163 63
163 37
3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
306 8 572 45
310 12 569 40
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 4
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
360 235 395 255
364 239 392 253
4 ____
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 130
44 278 580 322
48 282 576 314
130 MOD-8 synchronous up/down counter. The counter counts up when the 
control input = 1; it counts down when the control input = 0.
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
