CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 10 100 9
4 70 635 395
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 393 635 502
25165842 0
0
6 Title:
5 Name:
0
0
0
5
5 SCOPE
12 185 111 0 1 11
0 6
0
0 0 57584 0
1 D
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SCOPE
12 223 111 0 1 11
0 2
0
0 0 57584 0
2 CP
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 312 111 0 1 11
0 7
0
0 0 57584 0
1 Q
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
12 D Flip-Flop~
219 271 175 0 4 9
0 6 2 9 7
0
0 0 4208 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6153 0 0
0
0
9 Data Seq~
170 119 123 0 17 18
0 10 11 12 13 14 15 6 2 16
17 1 1 51 10 11 0 52
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
5394 0 0
0
0
AAAAABAAACADACAAABAAACADACACADACAAABAAAAABACACADACACADACACADACACADACACADACACADAC
ACADACACADACACADACACADAC
10
8 2 2 0 0 12432 0 5 4 0 0 6
151 159
163 159
163 169
237 169
237 157
247 157
0 0 1 0 0 4272 0 0 0 0 0 2
454 114
454 164
0 0 3 0 0 4240 0 0 0 0 0 2
404 164
476 164
0 0 4 0 0 4240 0 0 0 0 0 2
404 130
476 130
0 0 5 0 0 4240 0 0 0 0 0 2
404 114
476 114
1 0 2 0 0 16 0 2 0 0 1 2
223 123
223 169
1 0 6 0 0 4112 0 1 0 0 8 2
185 123
185 139
7 1 6 0 0 12432 0 5 4 0 0 4
151 150
163 150
163 139
247 139
1 4 7 0 0 8336 0 3 4 0 0 3
312 123
312 139
295 139
0 0 8 0 0 4224 0 0 0 0 0 5
307 242
579 242
579 274
307 274
307 242
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 64
20 238 276 282
24 242 272 274
64 D Flip-flop that triggers only 
on positive-going transitions.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 28
402 111 482 175
406 115 478 163
28 D  CP  Q
0      0
1      1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
431 127 447 151
435 131 443 147
1 ^
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
431 125 447 149
435 129 443 145
1 |
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
431 144 447 168
435 148 443 164
1 ^
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
431 142 447 166
435 146 443 162
1 |
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
309 239 575 276
313 243 572 271
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 4.6e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
