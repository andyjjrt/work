CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 436 635 605
27262994 0
0
6 Title:
5 Name:
0
0
0
21
10 2-In NAND~
219 111 215 0 3 22
0 2 4 6
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
8953 0 0
0
0
2 +V
167 191 119 0 1 3
0 10
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
2 +V
167 288 118 0 1 3
0 9
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
2 +V
167 377 118 0 1 3
0 11
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
2 +V
167 468 118 0 1 3
0 12
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
5 SCOPE
12 491 70 0 1 11
0 8
0
0 0 57584 0
2 CP
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 397 70 0 1 11
0 7
0
0 0 57584 0
1 A
-4 -4 3 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 308 70 0 1 11
0 4
0
0 0 57584 0
1 B
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 216 70 0 1 11
0 3
0
0 0 57584 0
1 C
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 127 70 0 1 11
0 2
0
0 0 57584 0
1 D
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
5 SCOPE
12 209 203 0 1 11
0 6
0
0 0 57584 0
3 CLR
-11 -4 10 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
7 Pulser~
4 522 177 0 10 12
0 13 14 8 15 0 0 20 20 21
7
0
0 0 4144 512
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8903 0 0
0
0
14 Logic Display~
6 150 64 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 239 64 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 331 64 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 420 64 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
6 74112~
219 430 195 0 7 32
0 12 12 8 12 6 16 7
0
0 0 4208 512
7 74LS112
-3 -60 46 -52
3 U1A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 4 0
1 U
3874 0 0
0
0
6 74112~
219 341 195 0 7 32
0 11 11 7 11 6 17 4
0
0 0 4208 512
7 74LS112
-3 -60 46 -52
3 U1B
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 2 4 0
1 U
6671 0 0
0
0
6 74112~
219 252 195 0 7 32
0 9 9 4 9 6 18 3
0
0 0 4208 512
7 74LS112
-3 -60 46 -52
3 U2A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 5 0
1 U
3789 0 0
0
0
6 74112~
219 159 195 0 7 32
0 10 10 3 10 6 19 2
0
0 0 4208 512
7 74LS112
-3 -60 46 -52
3 U2B
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 2 5 0
1 U
4871 0 0
0
0
12 Hex Display~
7 87 54 0 16 19
10 7 4 3 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3750 0 0
0
0
37
4 0 2 0 0 4096 0 21 0 0 8 2
78 78
78 112
3 0 3 0 0 8320 0 21 0 0 18 3
84 78
84 104
216 104
2 0 4 0 0 4096 0 21 0 0 7 2
90 78
90 97
0 0 5 0 0 4224 0 0 0 0 0 5
298 271
569 271
569 303
298 303
298 271
1 0 6 0 0 0 0 11 0 0 12 2
209 215
209 215
1 0 7 0 0 8320 0 21 0 0 20 3
96 78
96 90
397 90
2 0 4 0 0 12416 0 1 0 0 19 4
87 224
66 224
66 97
308 97
1 0 2 0 0 8320 0 1 0 0 17 4
87 206
78 206
78 112
127 112
5 0 6 0 0 4096 0 20 0 0 12 2
159 207
159 215
5 0 6 0 0 0 0 19 0 0 12 2
252 207
252 215
5 0 6 0 0 0 0 18 0 0 12 2
341 207
341 215
3 5 6 0 0 4224 0 1 17 0 0 3
138 215
430 215
430 207
1 0 2 0 0 0 0 13 0 0 17 2
150 82
127 82
1 0 3 0 0 0 0 14 0 0 18 2
239 82
216 82
1 0 4 0 0 0 0 15 0 0 19 2
331 82
308 82
1 0 7 0 0 0 0 16 0 0 20 2
420 82
397 82
1 7 2 0 0 0 0 10 20 0 0 3
127 82
127 159
135 159
1 0 3 0 0 0 0 9 0 0 35 2
216 82
216 159
1 0 4 0 0 0 0 8 0 0 36 2
308 82
308 159
1 0 7 0 0 0 0 7 0 0 37 2
397 82
397 159
1 0 8 0 0 4224 0 6 0 0 22 2
491 82
491 168
3 3 8 0 0 0 0 12 17 0 0 2
498 168
460 168
2 0 9 0 0 4096 0 19 0 0 28 2
276 159
288 159
1 0 10 0 0 4096 0 20 0 0 26 2
159 132
191 132
2 0 10 0 0 0 0 20 0 0 26 2
183 159
191 159
4 1 10 0 0 8320 0 20 2 0 0 3
183 177
191 177
191 128
1 0 9 0 0 4096 0 19 0 0 28 2
252 132
288 132
4 1 9 0 0 8320 0 19 3 0 0 3
276 177
288 177
288 127
1 0 11 0 0 4096 0 18 0 0 31 2
341 132
377 132
2 0 11 0 0 0 0 18 0 0 31 2
365 159
377 159
1 4 11 0 0 4224 0 4 18 0 0 3
377 127
377 177
365 177
1 0 12 0 0 4096 0 17 0 0 34 2
430 132
468 132
2 0 12 0 0 0 0 17 0 0 34 2
454 159
468 159
1 4 12 0 0 4224 0 5 17 0 0 3
468 127
468 177
454 177
7 3 3 0 0 0 0 19 20 0 0 4
228 159
207 159
207 168
189 168
7 3 4 0 0 0 0 18 19 0 0 4
317 159
298 159
298 168
282 168
7 3 7 0 0 0 0 17 18 0 0 4
406 159
386 159
386 168
371 168
2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 31
15 278 271 302
19 282 267 298
31 MOD-10 (decade) ripple counter.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
300 268 566 305
304 272 563 300
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0159882 0 4.98503e-315 0 0.016 0.016
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
