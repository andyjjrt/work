CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 355
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 355 635 464
25165842 0
0
6 Title:
5 Name:
0
0
0
5
5 SCOPE
12 238 98 0 1 11
0 3
0
0 0 57568 0
1 A
-4 -4 3 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SCOPE
12 280 98 0 1 11
0 2
0
0 0 57568 0
1 B
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 370 97 0 1 11
0 4
0
0 0 57568 0
3 Out
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
9 Data Seq~
170 179 88 0 17 18
0 6 7 8 9 10 11 2 3 12
13 1 1 20 10 1 0 33
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
6153 0 0
0
0
AAAAAAABADACAAABADACAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
8 2-In OR~
219 313 133 0 3 22
0 3 2 4
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5394 0 0
0
0
6
1 0 2 0 0 4096 0 2 0 0 3 2
280 110
280 115
1 0 3 0 0 4096 0 1 0 0 4 2
238 110
238 124
7 2 2 0 0 4224 0 4 5 0 0 4
211 115
280 115
280 142
300 142
1 8 3 0 0 4224 0 5 4 0 0 2
300 124
211 124
1 3 4 0 0 4224 0 3 5 0 0 3
370 109
370 133
346 133
0 0 5 0 0 4224 0 0 0 0 0 5
289 193
558 193
558 224
289 224
289 193
3
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 16
15 204 151 228
19 208 147 224
16 2-input OR gate.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
291 190 557 227
295 194 554 222
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
356 133 444 157
360 137 440 153
10 Output=A+B
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 2e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
