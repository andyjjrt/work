CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 564
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 564
8388626 0
0
6 Title:
5 Name:
0
0
0
20
13 Logic Switch~
5 111 352 0 1 11
0 4
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
1 D
-27 -4 -20 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 111 334 0 1 11
0 3
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
1 A
-26 -3 -19 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 111 294 0 1 11
0 8
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
1 C
-26 -4 -19 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 111 276 0 1 11
0 9
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
1 B
-26 -5 -19 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 128 38 0 1 11
0 12
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-25 -5 -18 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 128 58 0 1 11
0 14
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 B
-25 -4 -18 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 128 86 0 1 11
0 13
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 C
-25 -3 -18 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 128 112 0 1 11
0 11
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
1 D
-24 -5 -17 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
14 Logic Display~
6 458 286 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
8 2-In OR~
219 382 315 0 3 22
0 5 6 2
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
7931 0 0
0
0
9 2-In NOR~
219 176 343 0 3 22
0 3 4 6
0
0 0 112 0
6 74LS02
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
9325 0 0
0
0
10 2-In XNOR~
219 176 285 0 3 22
0 9 8 7
0
0 0 112 0
4 4077
-7 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 589837
65 0 0 0 4 1 7 0
1 U
8903 0 0
0
0
9 3-In AND~
219 285 294 0 4 22
0 7 3 4 5
0
0 0 112 0
6 74LS11
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 6 0
1 U
3834 0 0
0
0
14 Logic Display~
6 455 52 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
9 Inverter~
13 210 58 0 2 22
0 14 19
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
7668 0 0
0
0
9 Inverter~
13 210 86 0 2 22
0 13 18
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
4718 0 0
0
0
9 4-In AND~
219 282 71 0 5 22
0 12 19 18 11 17
0
0 0 112 0
6 74LS21
-21 -28 21 -20
3 U1A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0
65 0 0 0 2 1 3 0
1 U
3874 0 0
0
0
9 4-In AND~
219 282 125 0 5 22
0 11 13 14 12 15
0
0 0 112 0
6 74LS21
-21 -28 21 -20
3 U1B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0
65 0 0 0 2 2 3 0
1 U
6671 0 0
0
0
9 2-In NOR~
219 273 170 0 3 22
0 12 11 16
0
0 0 112 0
6 74LS02
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3789 0 0
0
0
8 3-In OR~
219 370 80 0 4 22
0 17 15 16 10
0
0 0 112 0
4 4075
-14 -24 14 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 5 0
1 U
4871 0 0
0
0
26
3 1 2 0 0 4224 0 10 9 0 0 3
415 315
458 315
458 304
2 0 3 0 0 12416 0 13 0 0 8 5
261 294
219 294
219 307
139 307
139 334
3 0 4 0 0 12416 0 13 0 0 7 5
261 303
228 303
228 317
149 317
149 352
4 1 5 0 0 4224 0 13 10 0 0 4
306 294
361 294
361 306
369 306
3 2 6 0 0 4224 0 11 10 0 0 4
215 343
361 343
361 324
369 324
3 1 7 0 0 4224 0 12 13 0 0 2
215 285
261 285
1 2 4 0 0 0 0 1 11 0 0 2
123 352
163 352
1 1 3 0 0 0 0 2 11 0 0 2
123 334
163 334
1 2 8 0 0 4224 0 3 12 0 0 2
123 294
160 294
1 1 9 0 0 4224 0 4 12 0 0 2
123 276
160 276
1 4 10 0 0 8320 0 14 20 0 0 3
455 70
455 80
403 80
2 0 11 0 0 4096 0 19 0 0 23 3
260 179
162 179
162 112
1 0 12 0 0 8192 0 19 0 0 16 3
260 161
250 161
250 139
2 0 13 0 0 4224 0 18 0 0 24 3
258 121
184 121
184 86
3 0 14 0 0 4224 0 18 0 0 25 3
258 130
177 130
177 58
4 0 12 0 0 8192 0 18 0 0 26 3
258 139
169 139
169 38
5 2 15 0 0 8320 0 18 20 0 0 4
303 125
339 125
339 80
358 80
3 3 16 0 0 8320 0 19 20 0 0 4
312 170
348 170
348 89
357 89
5 1 17 0 0 4224 0 17 20 0 0 2
303 71
357 71
4 0 11 0 0 0 0 17 0 0 23 3
258 85
250 85
250 112
3 2 18 0 0 4224 0 17 16 0 0 4
258 76
239 76
239 86
231 86
2 2 19 0 0 4224 0 17 15 0 0 4
258 67
239 67
239 58
231 58
1 1 11 0 0 4224 0 8 18 0 0 2
140 112
258 112
1 1 13 0 0 0 0 7 16 0 0 2
140 86
195 86
1 1 14 0 0 0 0 6 15 0 0 2
140 58
195 58
1 1 12 0 0 4224 0 5 17 0 0 4
140 38
250 38
250 58
258 58
30
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
461 319 477 343
465 323 473 339
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
503 80 519 104
507 84 515 100
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
495 80 511 104
499 84 507 100
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
431 80 447 104
435 84 443 100
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
423 80 439 104
427 84 435 100
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
321 144 337 168
325 148 333 164
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
313 144 329 168
317 148 325 164
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
321 44 337 68
325 48 333 64
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
313 44 329 68
317 48 325 64
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
312 151 336 175
316 155 332 171
2 AD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
299 106 339 130
303 110 335 126
4 ABCD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
399 88 519 112
403 92 515 108
14 z=ABCD+ABCD+AD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
305 52 345 76
309 56 341 72
4 ABCD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
262 365 294 389
266 369 290 385
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
493 312 509 336
497 316 505 332
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
501 312 517 336
505 316 513 332
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
453 305 485 329
457 309 481 325
3 ___
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
413 319 517 343
417 323 513 339
12 z=AD(B+C)+AD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
289 317 305 341
293 321 301 337
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
281 317 297 341
285 321 293 337
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
249 310 281 334
253 314 277 330
3 ___
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
326 261 358 285
330 265 354 281
3 ___
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
221 252 253 276
225 256 249 272
3 ___
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
221 266 253 290
225 270 249 286
3 B+C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
302 275 366 299
306 279 362 295
7 AD(B+C)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
334 275 350 299
338 279 346 295
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
229 266 245 290
233 270 241 286
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
249 324 305 348
253 328 301 344
6 A+D=AD
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
259 191 291 215
263 195 287 211
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 67
37 416 581 440
41 420 577 436
67 Example showing how an XNOR gate may be used to simplify a circuit.
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
5.01587e-315 0 5.45005e-315 0 5.01587e-315 5.45005e-315
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
4.89465e-315 4.81264e-315 5.35472e-315 5.29283e-315 4.91275e-315 4.91275e-315
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
