CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 393
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 393
8388626 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 77 126 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21616 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
5 CLEAR
-54 -5 -19 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 77 42 0 1 11
0 5
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
3 SET
-39 -4 -18 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
5 4001~
219 135 117 0 3 22
0 2 4 3
0
0 0 112 0
4 4001
-14 -24 14 -16
3 U1B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
3618 0 0
0
0
5 4001~
219 135 51 0 3 22
0 5 3 2
0
0 0 112 0
4 4001
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
6153 0 0
0
0
14 Logic Display~
6 224 92 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 224 27 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
13 SR Flip-Flop~
219 414 243 0 4 9
0 9 10 11 12
0
0 0 4208 0
4 SRFF
-14 -53 14 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
10
0 1 2 0 0 8336 0 0 3 4 0 5
178 51
178 72
118 72
118 108
122 108
2 0 3 0 0 12432 0 4 0 0 3 5
122 60
104 60
104 93
179 93
179 117
1 3 3 0 0 16 0 5 3 0 0 3
224 110
224 117
174 117
1 3 2 0 0 16 0 6 4 0 0 3
224 45
224 51
174 51
2 1 4 0 0 4240 0 3 1 0 0 2
122 126
89 126
1 1 5 0 0 4240 0 4 2 0 0 2
122 42
89 42
0 0 1 0 0 4272 0 0 0 0 0 2
422 30
422 112
0 0 6 0 0 4240 0 0 0 0 0 2
332 112
504 112
0 0 7 0 0 4240 0 0 0 0 0 2
332 45
504 45
0 0 8 0 0 4240 0 0 0 0 0 2
332 30
504 30
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 119
331 26 515 170
335 30 511 142
119 Set  Clear   Output
 0     0    No change
 1     0     Q=1
 0     1     Q=0
 1     1    Invalid*

*produces Q=Q=0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
397 145 429 169
401 149 425 165
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
125 145 157 169
129 149 153 165
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
227 38 243 62
231 42 239 58
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
227 30 243 54
231 34 239 50
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
229 103 245 127
233 107 241 123
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
427 114 443 138
431 118 439 134
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
399 241 431 265
403 245 427 261
3 (c)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 64
38 201 270 265
42 205 266 253
64 (a) NOR gate latch
(b) truth table
(c) simplified block symbol
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 2e-005 1e-008 1e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
