CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 432 635 559
25165842 0
0
6 Title:
5 Name:
0
0
0
9
7 Pulser~
4 360 108 0 10 12
0 9 10 7 11 0 0 5 5 6
7
0
0 0 4640 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8953 0 0
0
0
2 +V
167 438 47 0 1 3
0 8
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
5 SCOPE
12 179 72 0 1 11
0 4
0
0 0 57568 0
3 CPa
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 272 72 0 1 11
0 3
0
0 0 57568 0
2 Qa
-7 -4 7 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
5 SCOPE
12 405 72 0 1 11
0 7
0
0 0 57568 0
3 CPb
-11 -4 10 4
2 U1
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 522 72 0 1 11
0 6
0
0 0 57568 0
2 Qb
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
6 74113~
219 474 107 0 6 22
0 8 7 8 8 12 6
0
0 0 4192 0
6 74F113
-22 -42 20 -34
3 U2A
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 5 0
1 U
9914 0 0
0
0
9 Data Seq~
170 113 81 0 17 18
0 13 14 15 16 17 18 5 4 19
20 1 1 32 5 6 0 33
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
3747 0 0
0
0
AAAAABACADAEAFAGAHAIAJAKALAMANAOAPBABBBCBDBEBFBGBHBIBJBKBLBMBNBOBP
12 D Flip-Flop~
219 227 135 0 4 9
0 5 4 21 3
0
0 0 4192 0
3 DFF
-10 -53 11 -45
2 U6
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
13
0 0 0 0 0 16 0 0 0 0 0 4
525 147
536 147
536 153
548 153
0 0 0 0 0 0 0 0 0 0 0 4
251 154
260 154
260 148
270 148
0 0 2 0 0 0 0 0 0 0 0 5
326 270
595 270
595 301
326 301
326 270
1 4 3 0 0 8320 0 4 9 0 0 3
272 84
272 99
251 99
1 0 4 0 0 4096 0 3 0 0 7 2
179 84
179 117
7 1 5 0 0 4224 0 8 9 0 0 4
145 108
196 108
196 99
203 99
8 2 4 0 0 4224 0 8 9 0 0 2
145 117
203 117
1 6 6 0 0 8320 0 6 7 0 0 3
522 84
522 90
498 90
1 0 7 0 0 4096 0 5 0 0 10 2
405 84
405 99
2 3 7 0 0 4224 0 7 1 0 0 2
443 99
384 99
4 0 8 0 0 4096 0 7 0 0 13 2
474 63
438 63
1 0 8 0 0 0 0 7 0 0 13 2
450 90
438 90
1 3 8 0 0 4224 0 2 7 0 0 3
438 56
438 108
450 108
6
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
328 267 594 304
332 271 591 299
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 173
8 228 304 332
12 232 300 312
173 Clocked FFs have a clock input (CP) 
that is active on either (a) the 
PGT or (b) the NGT.  The control 
inputs determine the effect of the 
active clock transition.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
161 160 193 184
165 164 189 180
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
416 160 448 184
420 164 444 180
3 (b)
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 25
337 139 519 159
341 143 516 157
25 CP is activated by an NGT
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 22
87 140 248 160
91 144 245 158
22 CP is activated by PGT
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
