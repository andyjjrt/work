CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 432
8388626 0
0
6 Title:
5 Name:
0
0
0
5
13 Logic Switch~
5 317 151 0 1 11
0 6
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 C
-22 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 317 114 0 1 11
0 5
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 B
-22 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 317 77 0 1 11
0 7
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-22 -1 -15 7
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
5 4073~
219 399 114 0 4 22
0 7 5 6 8
0
0 0 112 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 2 0
1 U
6153 0 0
0
0
14 Logic Display~
6 458 95 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
8
0 0 1 0 0 4256 0 0 0 4 2 2
179 44
179 190
0 0 2 0 0 4224 0 0 0 0 0 2
88 190
230 190
0 0 3 0 0 4224 0 0 0 0 0 2
88 61
230 61
0 0 4 0 0 4224 0 0 0 0 0 2
88 44
229 44
2 1 5 0 0 4224 0 4 2 0 0 2
375 114
329 114
3 1 6 0 0 8320 0 4 1 0 0 4
375 123
354 123
354 151
329 151
1 1 7 0 0 8336 0 4 3 0 0 4
375 105
354 105
354 77
329 77
1 4 8 0 0 8320 0 5 4 0 0 3
458 113
458 114
420 114
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 153
87 41 231 225
91 45 227 189
153 A   B   C   x=ABC
0   0   0     0
0   0   1     0
0   1   0     0
0   1   1     0
1   0   0     0
1   0   1     0
1   1   0     0
1   1   1     1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 50
99 248 507 272
103 252 503 268
50 Truth table and symbol for a three-input AND gate.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
433 117 481 141
437 121 477 137
5 x=ABC
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
