CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 436 635 583
27262994 0
0
6 Title:
5 Name:
0
0
0
18
14 Logic Display~
6 384 62 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8953 0 0
0
0
14 Logic Display~
6 295 62 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 203 62 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 114 62 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
7 Pulser~
4 486 168 0 10 12
0 12 13 6 14 0 0 20 20 21
7
0
0 0 4128 512
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5394 0 0
0
0
5 SCOPE
12 455 68 0 1 11
0 6
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 361 68 0 1 11
0 5
0
0 0 57568 0
1 A
-4 -4 3 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 272 68 0 1 11
0 4
0
0 0 57568 0
1 B
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 180 68 0 1 11
0 3
0
0 0 57568 0
1 C
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 91 68 0 1 11
0 2
0
0 0 57568 0
1 D
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
2 +V
167 432 109 0 1 3
0 10
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
2 +V
167 341 109 0 1 3
0 9
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
2 +V
167 252 109 0 1 3
0 7
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
0
0
2 +V
167 155 109 0 1 3
0 8
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
6 74113~
219 124 167 0 6 22
0 8 3 8 8 15 2
0
0 0 4704 512
7 74LS113
-25 -42 24 -34
3 U2B
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 2 2 0
1 U
7668 0 0
0
0
6 74113~
219 217 167 0 6 22
0 7 4 7 7 16 3
0
0 0 4704 512
7 74LS113
-25 -42 24 -34
3 U2A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 2 0
1 U
4718 0 0
0
0
6 74113~
219 395 167 0 6 22
0 10 6 10 10 17 5
0
0 0 4704 512
7 74LS113
-25 -42 24 -34
3 U1B
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 2 1 0
1 U
3874 0 0
0
0
6 74113~
219 306 167 0 6 22
0 9 5 9 9 18 4
0
0 0 4704 512
7 74LS113
-25 -42 24 -34
3 U1A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 1 0
1 U
6671 0 0
0
0
26
0 0 11 0 0 16 0 0 0 0 0 5
285 269
556 269
556 301
285 301
285 269
1 0 2 0 0 4096 0 4 0 0 6 2
114 80
91 80
1 0 3 0 0 4096 0 3 0 0 7 2
203 80
180 80
1 0 4 0 0 4096 0 2 0 0 8 2
295 80
272 80
1 0 5 0 0 4096 0 1 0 0 9 2
384 80
361 80
1 6 2 0 0 4224 0 10 15 0 0 3
91 80
91 150
98 150
1 0 3 0 0 4224 0 9 0 0 24 2
180 80
180 150
1 0 4 0 0 4224 0 8 0 0 25 2
272 80
272 150
1 0 5 0 0 4224 0 7 0 0 26 2
361 80
361 150
1 0 6 0 0 4224 0 6 0 0 11 2
455 80
455 159
3 2 6 0 0 0 0 5 17 0 0 2
462 159
424 159
1 0 7 0 0 4096 0 16 0 0 17 2
239 150
252 150
4 0 8 0 0 4096 0 15 0 0 15 2
122 123
155 123
1 0 8 0 0 0 0 15 0 0 15 2
146 150
155 150
3 1 8 0 0 8320 0 15 14 0 0 3
146 168
155 168
155 118
4 0 7 0 0 4096 0 16 0 0 17 2
215 123
252 123
3 1 7 0 0 8320 0 16 13 0 0 3
239 168
252 168
252 118
4 0 9 0 0 4096 0 18 0 0 20 2
304 123
341 123
1 0 9 0 0 0 0 18 0 0 20 2
328 150
341 150
1 3 9 0 0 4224 0 12 18 0 0 3
341 118
341 168
328 168
4 0 10 0 0 4096 0 17 0 0 23 2
393 123
432 123
1 0 10 0 0 0 0 17 0 0 23 2
417 150
432 150
1 3 10 0 0 4224 0 11 17 0 0 3
432 118
432 168
417 168
6 2 3 0 0 0 0 16 15 0 0 4
191 150
171 150
171 159
153 159
6 2 4 0 0 0 0 18 16 0 0 4
280 150
262 150
262 159
246 159
6 2 5 0 0 0 0 17 18 0 0 4
369 150
350 150
350 159
335 159
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
287 266 553 303
291 270 550 298
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 42
35 260 219 304
39 264 215 296
42 Four-bit asynchronous 
(ripple) counter.
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
