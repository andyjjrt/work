CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 428
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 428
8388626 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 125 149 0 1 11
0 9
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
2 y0
-27 -3 -13 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 125 65 0 1 11
0 10
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
2 x1
-27 -4 -13 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 125 94 0 1 11
0 7
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
2 x0
-26 -4 -12 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 125 128 0 1 11
0 8
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
2 y1
-27 -3 -13 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
5 4081~
219 291 106 0 3 22
0 5 6 4
0
0 0 112 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 2 0
1 U
5394 0 0
0
0
10 2-In XNOR~
219 194 140 0 3 22
0 7 9 6
0
0 0 112 0
4 4077
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
7734 0 0
0
0
10 2-In XNOR~
219 194 74 0 3 22
0 10 8 5
0
0 0 112 0
4 4077
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
9914 0 0
0
0
14 Logic Display~
6 345 74 0 1 2
10 4
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
16
0 0 2 0 0 24704 0 0 0 0 0 8
94 116
89 116
89 139
83 139
83 140
89 140
89 164
96 164
0 0 3 0 0 24704 0 0 0 0 0 8
94 55
89 55
89 77
83 77
83 78
89 78
89 102
96 102
1 3 4 0 0 8320 0 8 5 0 0 3
345 92
345 106
312 106
1 3 5 0 0 8320 0 5 7 0 0 4
267 97
246 97
246 74
233 74
3 2 6 0 0 8320 0 6 5 0 0 4
233 140
246 140
246 115
267 115
1 1 7 0 0 8320 0 6 3 0 0 4
178 131
167 131
167 94
137 94
2 1 8 0 0 8320 0 7 4 0 0 4
178 83
145 83
145 128
137 128
2 1 9 0 0 4224 0 6 1 0 0 2
178 149
137 149
1 1 10 0 0 4224 0 7 2 0 0 2
178 65
137 65
0 0 11 0 0 4224 0 0 0 0 0 2
377 231
577 231
0 0 12 0 0 4224 0 0 0 0 0 2
377 166
577 166
0 0 13 0 0 4224 0 0 0 0 0 2
377 102
577 102
0 0 1 0 0 4256 0 0 0 0 0 2
501 22
501 297
0 0 14 0 0 4224 0 0 0 0 0 2
377 297
577 297
0 0 15 0 0 4224 0 0 0 0 0 2
377 22
577 22
0 0 16 0 0 4224 0 0 0 0 0 2
377 40
577 40
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 80
16 211 344 255
20 215 340 247
80 Circuit for detecting equality of two 
two-bit binary numbers and truth table.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 377
377 19 585 363
381 23 581 295
377 x1  x0  y1  y0  z(Output)
0   0   0   0      1
0   0   0   1      0
0   0   1   0      0
0   0   1   1      0
0   1   0   0      0
0   1   0   1      1
0   1   1   0      0
0   1   1   1      0
1   0   0   0      0
1   0   0   1      0
1   0   1   0      1
1   0   1   1      0
1   1   0   0      0
1   1   0   1      0
1   1   1   0      0
1   1   1   1      1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
17 120 81 164
21 124 77 156
14 Binary
number
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
17 58 81 102
21 62 77 94
14 Binary
number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
335 107 351 131
339 111 347 127
1 z
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 2e-005 1e-008 1e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
