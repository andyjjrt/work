CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 436
10485778 0
0
6 Title:
5 Name:
0
0
0
15
13 Logic Switch~
5 251 82 0 1 11
0 15
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
2 A3
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 251 97 0 1 11
0 14
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
2 A2
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 251 112 0 1 11
0 13
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
2 A1
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 251 127 0 1 11
0 12
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
2 A0
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 251 158 0 1 11
0 11
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
2 B3
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 251 173 0 1 11
0 10
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
2 B2
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 251 188 0 1 11
0 9
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
2 B1
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 251 204 0 1 11
0 3
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
2 B0
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
7 Ground~
168 310 217 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
4 4008
219 343 147 0 14 29
0 15 14 13 12 11 10 9 3 2
5 6 7 8 4
0
0 0 5216 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
16 4-bit Full Adder
-57 -94 55 -86
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 0 1 0 0 0
1 U
7931 0 0
0
0
14 Logic Display~
6 436 93 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
14 Logic Display~
6 453 93 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8903 0 0
0
0
14 Logic Display~
6 470 93 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 487 93 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3363 0 0
0
0
14 Logic Display~
6 402 93 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
14
1 9 2 0 0 4224 0 9 10 0 0 3
310 211
310 183
311 183
1 8 3 0 0 4224 0 8 10 0 0 4
263 204
301 204
301 174
311 174
1 14 4 0 0 4224 0 15 10 0 0 2
402 111
375 111
1 10 5 0 0 8320 0 14 10 0 0 3
487 111
487 156
375 156
1 11 6 0 0 8320 0 13 10 0 0 3
470 111
470 147
375 147
1 12 7 0 0 8320 0 12 10 0 0 3
453 111
453 138
375 138
1 13 8 0 0 8320 0 11 10 0 0 3
436 111
436 129
375 129
7 1 9 0 0 12416 0 10 7 0 0 4
311 165
291 165
291 188
263 188
6 1 10 0 0 4224 0 10 6 0 0 4
311 156
281 156
281 173
263 173
5 1 11 0 0 4224 0 10 5 0 0 4
311 147
272 147
272 158
263 158
4 1 12 0 0 4224 0 10 4 0 0 4
311 138
272 138
272 127
263 127
3 1 13 0 0 4224 0 10 3 0 0 4
311 129
280 129
280 112
263 112
2 1 14 0 0 12416 0 10 2 0 0 4
311 120
291 120
291 97
263 97
1 1 15 0 0 4224 0 1 10 0 0 4
263 82
301 82
301 111
311 111
4
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
243 287 347 311
247 291 343 307
12 4-bit adder.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 44
408 166 527 220
412 170 524 212
44 Sum appears at 
S3, S2, S1, S0 
outputs.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 30
78 158 214 202
82 162 210 194
30 Addend bits 
from B register
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 30
76 84 212 128
80 88 208 120
30 Augend bits 
from A register
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
