CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 473
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 473
8912918 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 48 195 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21616 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 A
-28 -3 -21 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 49 236 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21616 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 B
-29 -3 -22 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
12 NPN Trans:B~
219 162 195 0 3 7
0 9 10 8
0
0 0 592 0
6 2N2270
7 0 49 8
2 Q2
8 -1 22 7
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3618 0 0
0
0
12 NPN Trans:B~
219 214 162 0 3 7
0 12 9 11
0
0 0 592 0
6 2N2270
7 0 49 8
2 Q3
9 -2 23 6
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
6153 0 0
0
0
6 Diode~
219 219 194 0 2 5
0 11 3
0
0 0 592 270
5 DIODE
11 0 46 8
2 D1
12 -5 26 3
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
5394 0 0
0
0
12 NPN Trans:B~
219 214 238 0 3 7
0 3 8 2
0
0 0 592 0
6 2N2270
7 0 49 8
2 Q4
8 -3 22 5
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
7734 0 0
0
0
6 Diode~
219 83 195 0 2 5
0 7 6
0
0 0 592 180
5 DIODE
11 0 46 8
2 D2
-7 -18 7 -10
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
9914 0 0
0
0
2 +V
167 196 81 0 1 3
0 4
0
0 0 53616 0
3 +5V
-10 -15 11 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
7 Ground~
168 219 305 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
11 Multimeter~
205 283 173 0 21 21
0 3 21 22 2 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
7 Ground~
168 308 224 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
6 Diode~
219 83 236 0 2 5
0 7 5
0
0 0 592 180
5 DIODE
11 0 46 8
2 D3
-7 -18 7 -10
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
8903 0 0
0
0
6 Diode~
219 126 195 0 2 5
0 7 10
0
0 0 592 692
5 DIODE
11 0 46 8
2 D4
-7 -18 7 -10
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3834 0 0
0
0
9 Terminal~
194 275 213 0 1 3
0 3
0
0 0 49520 270
1 X
-7 -14 0 -6
2 T1
3 -17 17 -9
0
2 X;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
3363 0 0
0
0
9 Resistor~
219 104 123 0 3 5
0 4 7 1
0
0 0 880 270
2 4k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 167 121 0 3 5
0 4 9 1
0
0 0 880 270
4 1.6k
8 0 36 8
2 R2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 219 120 0 3 5
0 4 12 1
0
0 0 880 270
3 130
7 0 28 8
2 R4
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 167 267 0 4 5
0 8 2 0 -1
0
0 0 880 270
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
31
1 0 3 0 0 4096 0 10 0 0 2 2
258 196
258 212
0 1 3 0 0 4224 0 0 14 18 0 2
219 212
263 212
1 0 2 0 0 4096 0 9 0 0 10 2
219 299
219 293
1 0 4 0 0 4096 0 8 0 0 13 2
196 90
196 95
1 2 5 0 0 4224 0 2 12 0 0 2
61 236
73 236
2 1 6 0 0 4224 0 7 1 0 0 2
73 195
60 195
1 0 7 0 0 4096 0 13 0 0 9 2
116 195
104 195
1 0 7 0 0 0 0 7 0 0 9 2
93 195
104 195
2 1 7 0 0 4224 0 15 12 0 0 3
104 141
104 236
93 236
2 3 2 0 0 8320 0 18 6 0 0 4
167 285
167 293
219 293
219 256
1 4 2 0 0 16 0 11 10 0 0 2
308 218
308 196
1 0 4 0 0 4096 0 16 0 0 13 2
167 103
167 95
1 1 4 0 0 8320 0 15 17 0 0 4
104 105
104 95
219 95
219 102
2 0 8 0 0 4096 0 6 0 0 17 2
196 238
167 238
2 0 9 0 0 4096 0 4 0 0 21 2
196 162
167 162
2 2 10 0 0 4224 0 13 3 0 0 2
136 195
144 195
3 1 8 0 0 4224 0 3 18 0 0 2
167 213
167 249
2 1 3 0 0 0 0 5 6 0 0 2
219 204
219 220
3 1 11 0 0 4224 0 4 5 0 0 2
219 180
219 184
2 1 12 0 0 4224 0 17 4 0 0 2
219 138
219 144
2 1 9 0 0 4224 0 16 3 0 0 2
167 139
167 177
0 0 1 0 0 4128 0 0 0 24 27 2
471 28
471 140
0 0 1 0 0 4256 0 0 0 28 31 2
471 191
471 319
0 0 13 0 0 4224 0 0 0 0 0 2
335 28
590 28
0 0 14 0 0 4224 0 0 0 0 0 2
335 56
590 56
0 0 15 0 0 4224 0 0 0 0 0 2
335 98
590 98
0 0 16 0 0 4224 0 0 0 0 0 2
335 140
590 140
0 0 17 0 0 4224 0 0 0 0 0 2
336 191
591 191
0 0 18 0 0 4224 0 0 0 0 0 2
337 219
592 219
0 0 19 0 0 4224 0 0 0 0 0 2
337 261
592 261
0 0 20 0 0 4224 0 0 0 0 0 2
337 319
592 319
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 60
14 299 182 363
18 303 178 351
60 TTL NAND gate with 
(a) LOW output and 
(b) HIGH output.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
451 322 479 342
455 326 476 340
3 (b)
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
451 145 479 165
455 149 476 163
3 (a)
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 195
362 23 579 162
366 27 576 139
195     Input          Output
  conditions     conditions
 A and B are
  both HIGH        Q3 OFF
   (>= 2V)
Input currents    Q4 ON so
 are very low    that Vx is
  IIH = 10uA    LOW (<= 0.4V)
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 280
334 187 600 343
338 191 597 317
280       Input              Output
    conditions         conditions
  A or B or both
     are LOW             Q4 OFF
    (<= 0.8V)
Current flows back     Q3 acts as
to ground through   emitter-follower
LOW input terminal  and VOH >= 2.4V,
   IIL = 1.1mA       typically 3.6V
22 .OPTIONS RSHUNT=1E12

1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
270270842 1210432 100 100 0 0
77 66 587 156
8 92 169 162
587 66
77 66
587 66
587 156
0 0
0.006 0 5.4 0 0.006 5.4
12401 0
4 0.003 2
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 15 -15 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
