CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 100 9
4 70 635 455
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 455 635 583
25165842 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 171 54 0 1 11
0 7
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 S
-24 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 171 71 0 1 11
0 6
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 E
-24 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
7 74LS157
122 287 155 0 14 29
0 7 15 14 13 12 11 10 9 8
6 5 4 3 2
0
0 0 4448 0
8 74ALS157
-27 -60 29 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 1 0 0 0
1 U
3618 0 0
0
0
9 Data Seq~
170 186 155 0 17 18
0 15 14 13 12 11 10 9 8 17
18 29 1 256 5 2 0 257
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
6153 0 0
0
0
AAAAABACADAEAFAGAHAIAJAKALAMANAOAPBABBBCBDBEBFBGBHBIBJBKBLBMBNBOBPCACBCCCDCECFCG
CHCICJCKCLCMCNCOCPDADBDCDDDEDFDGDHDIDJDKDLDMDNDODPEAEBECEDEEEFEGEHEIEJEKELEMENEO
EPFAFBFCFDFEFFFGFHFIFJFKFLFMFNFOFPGAGBGCGDGEGFGGGHGIGJGKGLGMGNGOGPHAHBHCHDHEHFHG
HHHIHJHKHLHMHNHOHPIAIBICIDIEIFIGIHIIIJIKILIMINIOIPJAJBJCJDJEJFJGJHJIJJJKJLJMJNJO
JPKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPLALBLCLDLELFLGLHLILJLKLLLMLNLOLPMAMBMCMDMEMFMG
MHMIMJMKMLMMMNMOMPNANBNCNDNENFNGNHNINJNKNLNMNNNONPOAOBOCODOEOFOGOHOIOJOKOLOMONOO
OPPAPBPCPDPEPFPGPHPIPJPKPLPMPNPOPP
5 SCOPE
12 336 117 0 1 11
0 5
0
0 0 57568 0
2 Za
-8 -4 6 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 361 132 0 1 11
0 4
0
0 0 57568 0
2 Zb
-8 -4 6 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 385 147 0 1 11
0 3
0
0 0 57568 0
2 Zc
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 410 162 0 1 11
0 2
0
0 0 57568 0
2 Zd
-8 -4 6 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
15
0 0 16 0 0 16 0 0 0 0 0 5
312 288
583 288
583 320
312 320
312 288
1 14 2 0 0 8320 0 8 3 0 0 3
410 174
410 191
319 191
1 13 3 0 0 8320 0 7 3 0 0 3
385 159
385 173
319 173
1 12 4 0 0 8320 0 6 3 0 0 3
361 144
361 155
319 155
1 11 5 0 0 8320 0 5 3 0 0 3
336 129
336 137
319 137
1 10 6 0 0 8320 0 2 3 0 0 4
183 71
233 71
233 200
249 200
1 1 7 0 0 8320 0 1 3 0 0 4
183 54
241 54
241 119
255 119
8 9 8 0 0 4224 0 4 3 0 0 2
218 191
255 191
7 8 9 0 0 4224 0 4 3 0 0 2
218 182
255 182
6 7 10 0 0 4224 0 4 3 0 0 2
218 173
255 173
5 6 11 0 0 4224 0 4 3 0 0 2
218 164
255 164
4 5 12 0 0 4224 0 4 3 0 0 2
218 155
255 155
3 4 13 0 0 4224 0 4 3 0 0 2
218 146
255 146
2 3 14 0 0 4224 0 4 3 0 0 2
218 137
255 137
1 2 15 0 0 4224 0 4 3 0 0 2
218 128
255 128
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
314 285 580 322
318 289 577 317
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 25
25 285 233 309
29 289 229 305
25 Quad 2-input multiplexer.
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
267780172 8525888 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
9.98039 0 5.4 0 10 10
12401 0
4 1e-006 2
2
221 112
0 7 0 0 2	0 16 0 0
367 106
0 2 0 0 1	0 16 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 16 0 0
200 112
0 7 0 0 2	0 16 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
