CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 436 635 587
27262994 0
0
6 Title:
5 Name:
0
0
0
23
2 +V
167 196 22 0 1 3
0 8
0
0 0 53616 0
3 +5V
-11 -13 10 -5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
4 LED~
171 369 83 0 2 2
10 8 11
0
0 0 112 0
4 LED1
17 0 45 8
2 D3
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
4441 0 0
0
0
4 LED~
171 283 83 0 2 2
10 8 10
0
0 0 112 0
4 LED1
17 0 45 8
2 D2
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
3618 0 0
0
0
4 LED~
171 196 83 0 2 2
10 8 9
0
0 0 112 0
4 LED1
17 0 45 8
2 D1
24 -10 38 -2
0
0
11 %D %1 %2 %M
0
0
4 SIP2
5

0 1 2 1 2 0
68 0 0 0 1 0 0 0
1 D
6153 0 0
0
0
9 Inverter~
13 347 98 0 2 22
0 4 11
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U9C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
5394 0 0
0
0
9 Inverter~
13 259 98 0 2 22
0 5 10
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U9B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
7734 0 0
0
0
9 Inverter~
13 169 98 0 2 22
0 6 9
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U9A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
9914 0 0
0
0
7 Pulser~
4 462 152 0 10 12
0 15 16 3 17 0 0 20 20 21
7
0
0 0 4144 512
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3747 0 0
0
0
5 SCOPE
12 426 69 0 1 11
0 3
0
0 0 57584 0
2 CP
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 326 69 0 1 11
0 4
0
0 0 57584 0
1 A
-4 -4 3 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
5 SCOPE
12 237 69 0 1 11
0 5
0
0 0 57584 0
1 B
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
5 SCOPE
12 149 69 0 1 11
0 6
0
0 0 57584 0
1 C
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
5 SCOPE
12 323 179 0 1 11
0 7
0
0 0 57584 0
3 CLR
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
2 +V
167 403 93 0 1 3
0 14
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
2 +V
167 312 93 0 1 3
0 13
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
2 +V
167 223 93 0 1 3
0 12
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
6 74112~
219 365 170 0 7 32
0 14 14 3 14 7 18 4
0
0 0 4208 512
7 74LS112
-3 -60 46 -52
3 U1A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 1 0
1 U
3874 0 0
0
0
6 74112~
219 276 170 0 7 32
0 13 13 4 13 7 19 5
0
0 0 4208 512
7 74LS112
-3 -60 46 -52
3 U1B
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 2 1 0
1 U
6671 0 0
0
0
6 74112~
219 187 170 0 7 32
0 12 12 5 12 7 20 6
0
0 0 4208 512
7 74LS112
-3 -60 46 -52
3 U2A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 2 0
1 U
3789 0 0
0
0
10 2-In NAND~
219 144 191 0 3 22
0 6 5 7
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4871 0 0
0
0
13 ResistorWire~
94 369 56 0 3 5
0 8 8 1
13 ResistorWire~
1 0 4400 270
3 330
5 -5 26 3
2 R3
6 -5 20 3
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 0 1 0 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
13 ResistorWire~
94 283 56 0 3 5
0 8 8 1
13 ResistorWire~
2 0 4400 270
3 330
5 -5 26 3
2 R2
6 -5 20 3
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 0 1 0 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
13 ResistorWire~
94 196 56 0 3 5
0 8 8 1
13 ResistorWire~
3 0 4400 270
3 330
5 -5 26 3
2 R1
6 -5 20 3
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 0 1 0 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
35
0 0 2 0 0 4240 0 0 0 0 0 5
305 270
576 270
576 301
305 301
305 270
1 0 3 0 0 4224 0 9 0 0 24 2
426 81
426 143
1 0 4 0 0 4096 0 10 0 0 15 2
326 81
326 98
1 0 5 0 0 4096 0 11 0 0 16 2
237 81
237 98
1 0 6 0 0 4096 0 12 0 0 17 2
149 81
149 98
0 1 6 0 0 8320 0 0 20 17 0 4
149 134
113 134
113 182
120 182
0 2 5 0 0 8320 0 0 20 34 0 5
237 143
237 215
113 215
113 200
120 200
1 0 7 0 0 0 0 13 0 0 23 2
323 191
323 191
1 0 8 0 0 4096 0 22 0 0 10 2
283 38
283 34
0 1 8 0 0 4224 0 0 21 13 0 3
196 34
369 34
369 38
2 1 8 0 0 0 0 21 2 0 0 2
369 74
369 73
2 1 8 0 0 0 0 22 3 0 0 2
283 74
283 73
1 1 8 0 0 0 0 1 23 0 0 2
196 31
196 38
2 1 8 0 0 0 0 23 4 0 0 2
196 74
196 73
1 0 4 0 0 8320 0 5 0 0 35 3
332 98
326 98
326 134
1 0 5 0 0 0 0 6 0 0 34 3
244 98
237 98
237 134
1 7 6 0 0 0 0 7 19 0 0 4
154 98
149 98
149 134
163 134
2 2 9 0 0 4224 0 7 4 0 0 3
190 98
196 98
196 93
2 2 10 0 0 8320 0 6 3 0 0 3
280 98
283 98
283 93
2 2 11 0 0 8320 0 5 2 0 0 3
368 98
369 98
369 93
5 0 7 0 0 4096 0 19 0 0 23 2
187 182
187 191
5 0 7 0 0 0 0 18 0 0 23 2
276 182
276 191
3 5 7 0 0 4224 0 20 17 0 0 3
171 191
365 191
365 182
3 3 3 0 0 0 0 8 17 0 0 2
438 143
395 143
2 0 12 0 0 4096 0 19 0 0 27 2
211 134
223 134
1 0 12 0 0 4096 0 19 0 0 27 2
187 107
223 107
4 1 12 0 0 8320 0 19 16 0 0 3
211 152
223 152
223 102
1 0 13 0 0 4096 0 18 0 0 30 2
276 107
312 107
2 0 13 0 0 0 0 18 0 0 30 2
300 134
312 134
1 4 13 0 0 4224 0 15 18 0 0 3
312 102
312 152
300 152
1 0 14 0 0 4096 0 17 0 0 33 2
365 107
403 107
2 0 14 0 0 0 0 17 0 0 33 2
389 134
403 134
1 4 14 0 0 4224 0 14 17 0 0 3
403 102
403 152
389 152
7 3 5 0 0 0 0 18 19 0 0 4
252 134
237 134
237 143
217 143
7 3 4 0 0 0 0 17 18 0 0 4
341 134
326 134
326 143
306 143
2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 58
14 266 270 310
18 270 266 302
58 LEDs are often used to display 
the states of a counter.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
307 267 573 304
311 271 570 299
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
