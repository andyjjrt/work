CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 432
8388626 0
0
6 Title:
5 Name:
0
0
0
5
13 Logic Switch~
5 121 149 0 1 11
0 2
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 B
-22 -2 -15 6
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 121 168 0 1 11
0 4
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 C
-22 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 121 130 0 1 11
0 5
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-22 -1 -15 7
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
14 Logic Display~
6 250 131 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
8 3-In OR~
219 176 149 0 4 22
0 5 2 4 3
0
0 0 96 0
4 4075
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 2 0
1 U
5394 0 0
0
0
8
2 1 2 0 0 4224 0 5 1 0 0 2
164 149
133 149
1 4 3 0 0 4224 0 4 5 0 0 2
250 149
209 149
3 1 4 0 0 12416 0 5 2 0 0 4
163 158
149 158
149 168
133 168
1 1 5 0 0 12416 0 5 3 0 0 4
163 140
149 140
149 130
133 130
0 0 1 0 0 4256 0 0 0 8 6 2
417 69
417 216
0 0 6 0 0 4224 0 0 0 0 0 2
323 216
488 216
0 0 7 0 0 4224 0 0 0 0 0 2
488 86
323 86
0 0 8 0 0 4224 0 0 0 0 0 2
323 69
490 69
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 49
89 267 489 291
93 271 485 287
49 Symbol and truth table for a three-inout OR gate.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 55
421 66 485 250
425 70 481 214
55 x=A+B+C
   0
   1
   1
   1
   1
   1
   1
   1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
330 66 354 250
334 70 350 214
25 A
0
0
0
0
1
1
1
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
390 67 414 251
394 71 410 215
25 C
0
1
0
1
0
1
0
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
359 66 383 250
363 70 379 214
25 B
0
0
1
1
0
0
1
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
221 152 285 176
225 156 281 172
7 x=A+B+C
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
