CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 20 100 9
4 70 635 556
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 556 635 628
25165842 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 218 30 0 1 11
0 28
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
2 S3
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 218 80 0 1 11
0 25
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
2 S0
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 218 63 0 1 11
0 26
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
2 S1
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 218 47 0 1 11
0 27
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
2 S2
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
14 Logic Display~
6 518 229 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
5 SCOPE
12 495 235 0 1 11
0 3
0
0 0 57584 0
1 X
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
9 Data Seq~
170 233 301 0 17 18
0 19 18 17 16 15 14 13 12 29
30 1 1 256 5 6 0 257
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS2
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
9914 0 0
0
0
AAAAABACADAEAFAGAHAIAJAKALAMANAOAPBABBBCBDBEBFBGBHBIBJBKBLBMBNBOBPCACBCCCDCECFCG
CHCICJCKCLCMCNCOCPDADBDCDDDEDFDGDHDIDJDKDLDMDNDODPEAEBECEDEEEFEGEHEIEJEKELEMENEO
EPFAFBFCFDFEFFFGFHFIFJFKFLFMFNFOFPGAGBGCGDGEGFGGGHGIGJGKGLGMGNGOGPHAHBHCHDHEHFHG
HHHIHJHKHLHMHNHOHPIAIBICIDIEIFIGIHIIIJIKILIMINIOIPJAJBJCJDJEJFJGJHJIJJJKJLJMJNJO
JPKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPLALBLCLDLELFLGLHLILJLKLLLMLNLOLPMAMBMCMDMEMFMG
MHMIMJMKMLMMMNMOMPNANBNCNDNENFNGNHNINJNKNLNMNNNONPOAOBOCODOEOFOGOHOIOJOKOLOMONOO
OPPAPBPCPDPEPFPGPHPIPJPKPLPMPNPOPP
9 Data Seq~
170 231 164 0 17 18
0 4 5 6 7 8 9 10 11 31
32 1 1 256 5 6 0 257
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
3747 0 0
0
0
AAPPPOPNPMPLPKPJPIPHPGPFPEPDPCPBPAOPOOONOMOLOKOJOIOHOGOFOEODOCOBOANPNONNNMNLNKNJ
NINHNGNFNENDNCNBNAMPMOMNMMMLMKMJMIMHMGMFMEMDMCMBMALPLOLNLMLLLKLJLILHLGLFLELDLCLB
LAKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAJPJOJNJMJLJKJJJIJHJGJFJEJDJCJBJAIPIOINIMILIKIJ
IIIHIGIFIEIDICIBIAHPHOHNHMHLHKHJHIHHHGHFHEHDHCHBHAGPGOGNGMGLGKGJGIGHGGGFGEGDGCGB
GAFPFOFNFMFLFKFJFIFHFGFFFEFDFCFBFAEPEOENEMELEKEJEIEHEGEFEEEDECEBEADPDODNDMDLDKDJ
DIDHDGDFDEDDDCDBDACPCOCNCMCLCKCJCICHCGCFCECDCCCBCABPBOBNBMBLBKBJBIBHBGBFBEBDBCBB
BAAPAOANAMALAKAJAIAHAGAFAEADACABAA
7 74LS151
20 328 301 0 14 29
0 19 18 17 16 15 14 13 12 28
27 26 25 23 33
0
0 0 12528 0
7 74HC151
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
7 74LS151
20 327 164 0 14 29
0 4 5 6 7 8 9 10 11 22
27 26 25 24 34
0
0 0 12528 0
7 74HC151
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
8 2-In OR~
219 441 255 0 3 22
0 24 23 3
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9325 0 0
0
0
9 Inverter~
13 326 30 0 2 22
0 28 22
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8903 0 0
0
0
32
0 0 2 0 0 4224 0 0 0 0 0 5
315 391
586 391
586 424
315 424
315 391
1 0 3 0 0 8320 0 5 0 0 22 3
518 247
518 255
495 255
1 1 4 0 0 4224 0 8 10 0 0 2
263 137
295 137
2 2 5 0 0 4224 0 8 10 0 0 2
263 146
295 146
3 3 6 0 0 4224 0 8 10 0 0 2
263 155
295 155
4 4 7 0 0 4224 0 8 10 0 0 2
263 164
295 164
5 5 8 0 0 4224 0 8 10 0 0 2
263 173
295 173
6 6 9 0 0 4224 0 8 10 0 0 2
263 182
295 182
7 7 10 0 0 4224 0 8 10 0 0 2
263 191
295 191
8 8 11 0 0 4224 0 8 10 0 0 2
263 200
295 200
8 8 12 0 0 4224 0 7 9 0 0 2
265 337
296 337
7 7 13 0 0 4224 0 7 9 0 0 2
265 328
296 328
6 6 14 0 0 4224 0 7 9 0 0 2
265 319
296 319
5 5 15 0 0 4224 0 7 9 0 0 2
265 310
296 310
4 4 16 0 0 4224 0 7 9 0 0 2
265 301
296 301
3 3 17 0 0 4224 0 7 9 0 0 2
265 292
296 292
2 2 18 0 0 4224 0 7 9 0 0 2
265 283
296 283
1 1 19 0 0 4224 0 7 9 0 0 2
265 274
296 274
0 0 20 0 0 8320 0 0 0 0 0 8
172 22
167 22
167 55
161 55
161 56
167 56
167 88
174 88
0 0 21 0 0 24704 0 0 0 0 0 8
172 121
167 121
167 233
161 233
161 234
167 234
167 354
174 354
2 9 22 0 0 8320 0 12 10 0 0 4
347 30
369 30
369 137
365 137
1 3 3 0 0 0 0 6 11 0 0 3
495 247
495 255
474 255
13 2 23 0 0 8320 0 9 11 0 0 4
360 328
414 328
414 264
428 264
13 1 24 0 0 4224 0 10 11 0 0 4
359 191
414 191
414 246
428 246
12 0 25 0 0 4096 0 10 0 0 29 2
359 164
387 164
11 0 26 0 0 4096 0 10 0 0 30 2
359 155
381 155
10 0 27 0 0 4096 0 10 0 0 31 2
359 146
375 146
0 9 28 0 0 4224 0 0 9 32 0 5
290 30
290 225
369 225
369 274
366 274
1 12 25 0 0 8320 0 2 9 0 0 4
230 80
387 80
387 301
360 301
1 11 26 0 0 8320 0 3 9 0 0 4
230 63
381 63
381 292
360 292
1 10 27 0 0 8320 0 4 9 0 0 4
230 47
375 47
375 283
360 283
1 1 28 0 0 0 0 1 12 0 0 2
230 30
311 30
8
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 132
9 367 297 451
13 371 293 435
132 Two 74HC151s combined to form a 
16-input multiplexer. The output 
is determined by S3 which enables 
one of the multiplexers.
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
108 214 148 258
112 218 144 250
9 Data
 in
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
95 36 159 80
99 40 155 72
13 Input
select
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
263 333 284 353
267 337 281 351
2 I0
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
263 256 284 276
267 260 281 274
2 I7
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
259 196 280 216
263 200 277 214
2 I8
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
258 119 286 139
262 123 283 137
3 I15
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
317 388 583 425
321 392 580 420
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
267780172 8525888 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.0159882 0 5.36094e-315 0 0.016 0.016
12401 0
4 1e-006 2
2
221 112
0 7 0 0 2	0 33 0 0
367 106
0 2 0 0 1	0 33 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 33 0 0
200 112
0 7 0 0 2	0 33 0 0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
