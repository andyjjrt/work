CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 440
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 440 635 566
27262994 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 203 100 0 1 11
0 2
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
16 Debounced switch
-130 -4 -18 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
9 Inverter~
13 325 118 0 2 22
0 5 3
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
4441 0 0
0
0
5 SCOPE
12 266 128 0 1 11
0 5
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 284 73 0 1 11
0 2
0
0 0 57568 0
1 A
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
5 SCOPE
12 419 73 0 1 11
0 4
0
0 0 57568 0
1 Q
-4 -4 3 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 509 73 0 1 11
0 6
0
0 0 57568 0
1 X
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
7 Pulser~
4 213 158 0 10 12
0 8 9 5 10 0 0 5 5 6
7
0
0 0 4128 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9914 0 0
0
0
9 2-In AND~
219 464 109 0 3 22
0 4 5 6
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3747 0 0
0
0
12 D Flip-Flop~
219 373 136 0 4 9
0 2 3 11 4
0
0 0 4192 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
10
0 0 7 0 0 16 0 0 0 0 0 5
318 264
589 264
589 296
318 296
318 264
1 0 2 0 0 4096 0 4 0 0 10 2
284 85
284 100
2 2 3 0 0 4224 0 2 9 0 0 2
346 118
349 118
1 0 4 0 0 4096 0 5 0 0 9 2
419 85
419 100
1 0 5 0 0 4096 0 3 0 0 8 2
266 140
266 149
1 3 6 0 0 4224 0 6 8 0 0 3
509 85
509 109
485 109
0 1 5 0 0 4096 0 0 2 8 0 3
305 149
305 118
310 118
3 2 5 0 0 4224 0 7 8 0 0 4
237 149
432 149
432 118
440 118
4 1 4 0 0 4224 0 9 8 0 0 2
397 100
440 100
1 1 2 0 0 4224 0 1 9 0 0 2
215 100
349 100
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
320 261 586 298
324 265 583 293
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 4
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 116
21 245 293 329
25 249 289 313
116 An edge-triggered D flip-flop 
is used to synchronize the 
enabling of the AND gate to the 
NGTs of the clock.
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
