CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 8 100 9
4 70 635 393
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 393
8388626 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 187 91 0 1 11
0 8
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 B
-23 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
14 Logic Display~
6 320 131 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
5 4081~
219 276 158 0 3 22
0 9 12 10
0
0 0 112 0
4 4081
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
3618 0 0
0
0
5 4081~
219 276 100 0 3 22
0 8 9 11
0
0 0 112 0
4 4081
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
6153 0 0
0
0
7 Pulser~
4 142 137 0 10 12
0 13 14 9 15 0 0 5 5 6
7
0
0 0 4144 0
0
2 V4
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
5394 0 0
0
0
14 Logic Display~
6 320 74 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
9 Inverter~
13 226 167 0 2 22
0 8 12
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
9914 0 0
0
0
13
0 0 2 0 0 24704 0 0 0 0 0 8
388 135
383 135
383 151
377 151
377 152
383 152
383 169
390 169
0 0 3 0 0 20608 0 0 0 0 0 6
405 160
414 160
414 153
422 153
422 160
433 160
0 0 4 0 0 4224 0 0 0 0 0 2
405 142
433 142
0 0 5 0 0 24704 0 0 0 0 0 8
388 76
383 76
383 92
377 92
377 93
383 93
383 110
390 110
0 0 6 0 0 4224 0 0 0 0 0 2
405 101
433 101
0 0 7 0 0 20608 0 0 0 0 0 6
405 85
414 85
414 78
422 78
422 85
433 85
1 0 8 0 0 8320 0 7 0 0 8 3
211 167
200 167
200 91
1 1 8 0 0 0 0 4 1 0 0 2
252 91
199 91
3 0 9 0 0 4224 0 5 0 0 13 2
166 128
237 128
1 3 10 0 0 8320 0 2 3 0 0 3
320 149
320 158
297 158
3 1 11 0 0 4224 0 4 6 0 0 3
297 100
320 100
320 92
2 2 12 0 0 4224 0 3 7 0 0 2
252 167
247 167
2 1 9 0 0 0 0 4 3 0 0 4
252 109
237 109
237 149
252 149
12
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
392 149 406 169
396 153 403 167
1 0
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
392 131 406 151
396 135 403 149
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
434 145 490 169
438 149 486 165
6 IF B=0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
435 127 491 151
439 131 487 147
6 IF B=1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
392 90 406 110
396 94 403 108
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
434 86 490 110
438 90 486 106
6 IF B=0
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
392 74 406 94
396 78 403 92
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
434 70 490 94
438 74 486 90
6 IF B=1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 122
56 229 552 273
60 233 548 265
122 This circuit is called a pulse-steering circuit because it 
steers the input to one output or the other, depending on B.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
158 109 174 133
162 113 170 129
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
326 139 342 163
330 143 338 159
1 Y
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
326 81 342 105
330 85 338 101
1 X
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 2e-005 1e-008 1e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
