CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 436 635 587
27262994 0
0
6 Title:
5 Name:
0
0
0
16
14 Logic Display~
6 355 46 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8953 0 0
0
0
14 Logic Display~
6 266 46 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 174 46 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
7 Pulser~
4 462 152 0 10 12
0 11 12 6 13 0 0 20 20 21
7
0
0 0 4128 512
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6153 0 0
0
0
5 SCOPE
12 426 52 0 1 11
0 6
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 332 52 0 1 11
0 5
0
0 0 57568 0
1 A
-4 -4 3 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 243 52 0 1 11
0 4
0
0 0 57568 0
1 B
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 151 52 0 1 11
0 3
0
0 0 57568 0
1 C
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 235 180 0 1 11
0 2
0
0 0 57568 0
3 CLR
-11 -4 10 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
2 +V
167 403 93 0 1 3
0 9
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
2 +V
167 312 93 0 1 3
0 8
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
2 +V
167 223 93 0 1 3
0 7
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
6 74112~
219 365 170 0 7 32
0 9 9 6 9 2 14 5
0
0 0 4192 512
7 74LS112
-3 -60 46 -52
3 U1A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 1 0
1 U
3834 0 0
0
0
6 74112~
219 276 170 0 7 32
0 8 8 5 8 2 15 4
0
0 0 4192 512
7 74LS112
-3 -60 46 -52
3 U1B
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 2 1 0
1 U
3363 0 0
0
0
6 74112~
219 187 170 0 7 32
0 7 7 4 7 2 16 3
0
0 0 4192 512
7 74LS112
-3 -60 46 -52
3 U2A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 2 0
1 U
7668 0 0
0
0
10 2-In NAND~
219 144 191 0 3 22
0 4 3 2
0
0 0 608 0
6 74LS00
-14 -24 28 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4718 0 0
0
0
26
0 0 10 0 0 16 0 0 0 0 0 5
300 266
571 266
571 298
300 298
300 266
1 0 2 0 0 4096 0 9 0 0 7 2
235 192
235 191
0 2 3 0 0 8320 0 0 16 11 0 4
151 85
101 85
101 200
120 200
0 1 4 0 0 4224 0 0 16 12 0 4
243 75
112 75
112 182
120 182
5 0 2 0 0 4096 0 15 0 0 7 2
187 182
187 191
5 0 2 0 0 0 0 14 0 0 7 2
276 182
276 191
3 5 2 0 0 4224 0 16 13 0 0 3
171 191
365 191
365 182
1 0 3 0 0 0 0 3 0 0 11 2
174 64
151 64
1 0 4 0 0 0 0 2 0 0 12 2
266 64
243 64
1 0 5 0 0 4096 0 1 0 0 13 2
355 64
332 64
1 7 3 0 0 0 0 8 15 0 0 3
151 64
151 134
163 134
1 0 4 0 0 0 0 7 0 0 25 2
243 64
243 134
1 0 5 0 0 4224 0 6 0 0 26 2
332 64
332 134
1 0 6 0 0 4224 0 5 0 0 15 2
426 64
426 143
3 3 6 0 0 0 0 4 13 0 0 2
438 143
395 143
2 0 7 0 0 4096 0 15 0 0 18 2
211 134
223 134
1 0 7 0 0 4096 0 15 0 0 18 2
187 107
223 107
4 1 7 0 0 8320 0 15 12 0 0 3
211 152
223 152
223 102
1 0 8 0 0 4096 0 14 0 0 21 2
276 107
312 107
2 0 8 0 0 0 0 14 0 0 21 2
300 134
312 134
1 4 8 0 0 4224 0 11 14 0 0 3
312 102
312 152
300 152
1 0 9 0 0 4096 0 13 0 0 24 2
365 107
403 107
2 0 9 0 0 0 0 13 0 0 24 2
389 134
403 134
1 4 9 0 0 4224 0 10 13 0 0 3
403 102
403 152
389 152
7 3 4 0 0 0 0 14 15 0 0 4
252 134
233 134
233 143
217 143
7 3 5 0 0 0 0 13 14 0 0 4
341 134
321 134
321 143
306 143
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
302 263 568 300
306 267 565 295
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 90
19 251 275 315
23 255 271 303
90 MOD-6 counter produced by 
clearing a MOD-8 counter when 
a count of six (110) occurs.
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
