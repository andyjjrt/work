CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 432
8388626 0
0
6 Title:
5 Name:
0
0
0
3
13 Logic Switch~
5 304 138 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21616 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-24 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
14 Logic Display~
6 422 114 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
9 Inverter~
13 355 138 0 2 22
0 3 2
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 2 0
1 U
3618 0 0
0
0
6
2 1 2 0 0 4224 0 3 2 0 0 3
376 138
422 138
422 132
1 1 3 0 0 4224 0 1 3 0 0 2
316 138
340 138
0 0 1 0 0 4256 0 0 0 4 6 2
190 110
190 158
0 0 4 0 0 4224 0 0 0 0 0 2
159 110
222 110
0 0 5 0 0 4224 0 0 0 0 0 2
159 127
223 127
0 0 6 0 0 4224 0 0 0 0 0 2
159 158
223 158
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 60
124 258 476 302
128 262 472 294
60 (a) Truth table;
(b) symbol for the INVERTER (NOT circuit).
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
342 191 374 215
346 195 370 211
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
172 191 204 215
176 195 200 211
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
160 107 184 171
164 111 180 159
7 A
0
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
191 107 223 171
195 111 219 159
11 x=A
 1
 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
175 90 207 114
179 94 203 110
3 NOT
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
