CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 514
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 514
8388626 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 252 253 0 1 11
0 2
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
1 B
-23 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 252 235 0 1 11
0 3
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
1 A
-24 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 77 44 0 1 11
0 5
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-22 -5 -15 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 78 77 0 1 11
0 6
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 B
-23 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
14 Logic Display~
6 371 222 0 1 2
10 4
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
10 2-In XNOR~
219 299 244 0 3 22
0 3 2 4
0
0 0 112 0
4 4077
-7 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 589840
65 0 0 0 4 1 3 0
1 U
7734 0 0
0
0
5 4049~
219 152 77 0 2 22
0 6 7
0
0 0 112 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 2 2 0
1 U
9914 0 0
0
0
14 Logic Display~
6 333 54 0 1 2
10 14
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
9 2-In AND~
219 206 109 0 3 22
0 6 5 12
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3549 0 0
0
0
9 2-In AND~
219 206 53 0 3 22
0 11 7 13
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7931 0 0
0
0
5 4049~
219 151 44 0 2 22
0 5 11
0
0 0 112 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 2 0
1 U
9325 0 0
0
0
5 4071~
219 264 80 0 3 22
0 13 12 14
0
0 0 112 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 4 0
1 U
8903 0 0
0
0
16
2 1 2 0 0 4224 0 6 1 0 0 2
283 253
264 253
1 1 3 0 0 4224 0 6 2 0 0 2
283 235
264 235
1 3 4 0 0 8320 0 5 6 0 0 3
371 240
371 244
338 244
2 0 5 0 0 8320 0 9 0 0 12 3
182 118
112 118
112 44
1 0 6 0 0 4224 0 9 0 0 6 3
182 100
129 100
129 77
1 1 6 0 0 0 0 7 4 0 0 2
137 77
90 77
2 2 7 0 0 8320 0 10 7 0 0 3
182 62
173 62
173 77
0 0 1 0 0 4256 0 0 0 10 0 2
471 25
471 107
0 0 8 0 0 4224 0 0 0 0 0 2
413 107
494 107
0 0 9 0 0 4224 0 0 0 0 0 2
413 25
494 25
0 0 10 0 0 4224 0 0 0 0 0 2
413 41
492 41
1 1 5 0 0 0 0 11 3 0 0 2
136 44
89 44
1 2 11 0 0 4224 0 10 11 0 0 4
182 44
167 44
167 44
172 44
2 3 12 0 0 8320 0 12 9 0 0 4
251 89
232 89
232 109
227 109
1 3 13 0 0 4224 0 12 10 0 0 4
251 71
231 71
231 53
227 53
1 3 14 0 0 8320 0 8 12 0 0 3
333 72
333 80
297 80
27
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 81
84 350 428 394
88 354 424 386
81 (a) Exclusive-NOR circuit and truth table;
(b) traditional symbol for XNOR gate.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
477 21 501 125
481 25 497 105
13 x
1
0
0
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
444 21 468 125
448 25 464 105
13 B
0
1
0
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
417 21 441 125
421 25 437 105
13 A
0
0
1
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
238 44 254 68
242 48 250 64
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
348 77 364 101
352 81 360 97
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
340 77 356 101
344 81 352 97
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
300 85 364 109
304 89 360 105
7 x=AB+AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
230 52 254 76
234 56 250 72
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
230 90 254 114
234 94 250 110
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
230 44 246 68
234 48 242 64
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
174 35 190 59
178 39 186 55
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
174 17 190 41
178 21 186 37
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
173 25 189 49
177 29 185 45
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
174 43 190 67
178 47 186 63
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
174 100 190 124
178 104 186 120
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
175 81 191 105
179 85 187 101
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
294 119 326 143
298 123 322 139
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
296 287 328 311
300 291 324 307
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
363 255 379 279
367 259 375 275
1 +
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
363 255 379 279
367 259 375 275
1 O
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
345 269 401 293
349 273 397 289
6 =AB+AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
337 255 369 279
341 259 365 275
3 x=A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
374 255 390 279
378 259 386 275
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
385 261 401 285
389 265 397 281
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
352 240 392 264
356 244 388 260
4 ____
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
377 261 393 285
381 265 389 281
1 -
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
