CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 720 463
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 463 720 614
27262994 0
0
6 Title:
5 Name:
0
0
0
29
5 SCOPE
12 145 205 0 1 11
0 17
0
0 0 57584 0
2 CP
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
12 Hex Display~
7 34 45 0 16 19
10 5 4 3 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4441 0 0
0
0
14 Logic Display~
6 90 43 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 239 43 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
5 SCOPE
12 216 49 0 1 11
0 5
0
0 0 57584 0
1 A
-4 -4 3 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
14 Logic Display~
6 140 43 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
5 SCOPE
12 167 49 0 1 11
0 4
0
0 0 57584 0
1 B
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 117 49 0 1 11
0 3
0
0 0 57584 0
1 C
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 67 49 0 1 11
0 2
0
0 0 57584 0
1 D
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
14 Logic Display~
6 190 43 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
9 Terminal~
194 25 111 0 1 3
0 2
0
0 0 49520 180
1 D
-3 0 4 8
2 T1
3 -17 17 -9
0
2 D;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9325 0 0
0
0
9 Terminal~
194 31 111 0 1 3
0 3
0
0 0 49520 180
1 C
-3 0 4 8
2 T6
3 -17 17 -9
0
2 C;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8903 0 0
0
0
9 Terminal~
194 37 111 0 1 3
0 4
0
0 0 49520 180
1 B
-3 0 4 8
2 T7
3 -17 17 -9
0
2 B;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3834 0 0
0
0
9 Terminal~
194 43 111 0 1 3
0 5
0
0 0 49520 180
1 A
-3 0 4 8
2 T8
3 -17 17 -9
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3363 0 0
0
0
9 3-In AND~
219 265 83 0 4 22
0 5 4 3 18
0
0 0 112 512
6 74LS11
-21 -28 21 -20
3 U8A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 4 0
1 U
7668 0 0
0
0
9 2-In AND~
219 354 96 0 3 22
0 5 4 19
0
0 0 112 512
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4718 0 0
0
0
2 +V
167 203 143 0 1 3
0 20
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3874 0 0
0
0
6 74113~
219 205 191 0 6 22
0 18 17 18 20 24 2
0
0 0 4208 512
7 74LS113
-25 -42 24 -34
3 U2B
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 2 2 0
1 U
6671 0 0
0
0
6 74113~
219 295 190 0 6 22
0 19 17 19 21 25 3
0
0 0 4208 512
7 74LS113
-25 -42 24 -34
3 U2A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 2 0
1 U
3789 0 0
0
0
6 74113~
219 384 190 0 6 22
0 5 17 5 22 26 4
0
0 0 4208 512
7 74LS113
-25 -42 24 -34
3 U1B
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 2 1 0
1 U
4871 0 0
0
0
6 74113~
219 460 190 0 6 22
0 23 17 23 23 27 5
0
0 0 4208 512
7 74LS113
-25 -42 24 -34
3 U1A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 1 0
1 U
3750 0 0
0
0
2 +V
167 496 132 0 1 3
0 23
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8778 0 0
0
0
2 +V
167 382 143 0 1 3
0 22
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
538 0 0
0
0
2 +V
167 293 142 0 1 3
0 21
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6843 0 0
0
0
7 Pulser~
4 73 207 0 10 12
0 28 29 17 30 0 0 20 20 21
7
0
0 0 4144 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3136 0 0
0
0
9 Terminal~
194 429 165 0 1 3
0 5
0
0 0 49520 0
1 A
-4 -12 3 -4
2 T2
-7 -32 7 -24
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5950 0 0
0
0
9 Terminal~
194 351 165 0 1 3
0 4
0
0 0 49520 0
1 B
-3 -12 4 -4
2 T3
-7 -32 7 -24
0
2 B;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5670 0 0
0
0
9 Terminal~
194 261 165 0 1 3
0 3
0
0 0 49520 0
1 C
-3 -12 4 -4
2 T4
-7 -32 7 -24
0
2 C;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6828 0 0
0
0
9 Terminal~
194 174 165 0 1 3
0 2
0
0 0 49520 0
1 D
-3 -13 4 -5
2 T5
-7 -32 7 -24
0
2 D;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6735 0 0
0
0
50
0 0 6 0 0 4224 0 0 0 0 0 5
155 248
426 248
426 281
155 281
155 248
0 0 7 0 0 4224 0 0 0 0 0 2
658 11
658 340
0 0 8 0 0 4224 0 0 0 0 0 2
630 12
630 340
0 0 9 0 0 4224 0 0 0 0 0 2
595 12
595 340
0 0 1 0 0 4256 0 0 0 12 10 2
568 6
568 345
0 0 10 0 0 4224 0 0 0 0 0 2
515 278
683 278
0 0 11 0 0 4224 0 0 0 0 0 2
515 215
682 215
0 0 12 0 0 4224 0 0 0 0 0 2
515 150
682 150
0 0 13 0 0 4224 0 0 0 0 0 2
515 86
683 86
0 0 14 0 0 4224 0 0 0 0 0 2
515 345
682 345
0 0 15 0 0 4224 0 0 0 0 0 2
682 22
515 22
0 0 16 0 0 4224 0 0 0 0 0 2
515 6
684 6
1 0 17 0 0 4096 0 1 0 0 47 2
145 217
145 216
0 1 3 0 0 4224 0 0 8 19 0 3
31 84
117 84
117 61
0 1 4 0 0 4224 0 0 7 18 0 3
37 79
167 79
167 61
0 1 5 0 0 4224 0 0 5 17 0 3
43 74
216 74
216 61
1 1 5 0 0 0 0 2 14 0 0 2
43 69
43 96
2 1 4 0 0 0 0 2 13 0 0 2
37 69
37 96
3 1 3 0 0 0 0 2 12 0 0 2
31 69
31 96
4 1 2 0 0 4096 0 2 11 0 0 2
25 69
25 96
1 0 5 0 0 0 0 4 0 0 16 2
239 61
216 61
1 0 4 0 0 0 0 10 0 0 15 2
190 61
167 61
1 0 3 0 0 0 0 6 0 0 14 2
140 61
117 61
1 0 2 0 0 0 0 3 0 0 25 2
90 61
67 61
1 0 2 0 0 8320 0 9 0 0 20 3
67 61
67 89
25 89
1 6 2 0 0 0 0 29 18 0 0 2
174 174
179 174
1 0 3 0 0 0 0 28 0 0 30 2
261 174
261 173
1 0 4 0 0 0 0 27 0 0 37 2
351 174
351 173
1 0 5 0 0 0 0 26 0 0 40 2
429 174
429 173
3 6 3 0 0 0 0 15 19 0 0 6
285 92
290 92
290 124
252 124
252 173
269 173
2 0 4 0 0 0 0 15 0 0 37 4
285 83
314 83
314 124
342 124
1 0 5 0 0 0 0 15 0 0 38 3
285 74
387 74
387 87
4 0 18 0 0 8320 0 15 0 0 34 3
240 83
234 83
234 174
3 1 18 0 0 0 0 18 18 0 0 4
227 192
243 192
243 174
227 174
3 0 19 0 0 8320 0 16 0 0 36 3
329 96
323 96
323 173
3 1 19 0 0 0 0 19 19 0 0 4
317 191
332 191
332 173
317 173
2 6 4 0 0 0 0 16 20 0 0 5
374 105
374 124
342 124
342 173
358 173
1 0 5 0 0 0 0 16 0 0 40 3
374 87
420 87
420 173
3 0 5 0 0 0 0 20 0 0 40 3
406 191
420 191
420 173
1 6 5 0 0 0 0 20 21 0 0 2
406 173
434 173
1 4 20 0 0 4224 0 17 18 0 0 2
203 152
203 147
1 4 21 0 0 4224 0 24 19 0 0 2
293 151
293 146
1 4 22 0 0 4224 0 23 20 0 0 2
382 152
382 146
2 0 17 0 0 4096 0 18 0 0 47 2
234 183
234 216
2 0 17 0 0 4096 0 19 0 0 47 2
324 182
324 216
2 0 17 0 0 0 0 20 0 0 47 2
413 182
413 216
3 2 17 0 0 12416 0 25 21 0 0 5
97 198
114 198
114 216
489 216
489 182
4 0 23 0 0 4096 0 21 0 0 50 2
458 146
496 146
1 0 23 0 0 0 0 21 0 0 50 2
482 173
496 173
1 3 23 0 0 4224 0 22 21 0 0 3
496 141
496 191
482 191
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 105
517 3 565 427
521 7 561 343
105 Count
  0
  1
  2
  3
  4
  5
  6
  7
  8
  9
 10
 11
 12
 13
 14
 15
  0
  .
  .
  .
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 61
661 3 685 427
665 7 681 343
61 A
0
1
0
1
0
1
0
1
0
1
0
1
0
1
0
1
0
.
.
.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 61
636 3 660 427
640 7 656 343
61 B
0
0
1
1
0
0
1
1
0
0
1
1
0
0
1
1
0
.
.
.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 83
596 3 636 427
600 7 632 343
83  C
 0
 0
 0
 0
 1
 1
 1
 1
 0
 0
 0
 0
 1
 1
 1
 1
 0
 .
 .
etc
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 61
573 3 597 427
577 7 593 343
61 D
0
0
0
0
0
0
0
0
1
1
1
1
1
1
1
1
0
.
.
.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 134
5 294 493 358
9 298 489 346
134 Synchronous MOD-16 counter.  Each FF is clocked by the NGT 
of the clock input so that all FF transitions occur at the 
same time.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
157 245 423 282
161 249 420 277
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
