CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 440
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 440 635 591
27262994 0
0
6 Title:
5 Name:
0
0
0
22
9 Terminal~
194 330 161 0 1 3
0 2
0
0 0 49520 270
2 YN
-10 -13 4 -5
2 T6
-7 -25 7 -17
0
3 YN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8953 0 0
0
0
9 Terminal~
194 442 161 0 1 3
0 3
0
0 0 49520 270
2 ZN
-10 -13 4 -5
2 T5
-7 -25 7 -17
0
3 ZN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4441 0 0
0
0
9 Terminal~
194 292 241 0 1 3
0 3
0
0 0 49520 90
2 ZN
-20 -4 -6 4
2 T4
-7 -25 7 -17
0
3 ZN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3618 0 0
0
0
9 Terminal~
194 292 232 0 1 3
0 2
0
0 0 49520 90
2 YN
-20 -5 -6 3
2 T3
-7 -25 7 -17
0
3 YN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6153 0 0
0
0
9 Terminal~
194 218 143 0 1 3
0 4
0
0 0 49520 270
1 X
-7 -13 0 -5
2 T2
-7 -25 7 -17
0
2 X;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5394 0 0
0
0
9 Terminal~
194 292 223 0 1 3
0 4
0
0 0 49520 90
1 X
-14 -6 -7 2
2 T1
-7 -25 7 -17
0
2 X;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7734 0 0
0
0
5 SCOPE
12 216 193 0 1 11
0 8
0
0 0 57584 0
2 CP
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 4023~
219 327 230 0 4 22
0 4 2 3 5
0
0 0 112 0
4 4023
-14 -28 14 -20
3 U7A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 3 0
1 U
3747 0 0
0
0
14 Logic Display~
6 484 60 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 344 60 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7931 0 0
0
0
14 Logic Display~
6 224 60 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
6 74113~
219 178 159 0 6 22
0 10 7 10 10 13 4
0
0 0 4208 0
7 74LS113
-25 -42 24 -34
3 U1A
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 1 0
1 U
8903 0 0
0
0
6 74113~
219 288 159 0 6 22
0 9 6 9 9 2 7
0
0 0 4208 0
7 74LS113
-25 -42 24 -34
3 U1B
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 2 1 0
1 U
3834 0 0
0
0
6 74113~
219 401 159 0 6 22
0 5 8 5 11 3 6
0
0 0 4208 0
7 74LS113
-25 -42 24 -34
3 U2A
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 1 2 0
1 U
3363 0 0
0
0
2 +V
167 140 104 0 1 3
0 10
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
2 +V
167 249 104 0 1 3
0 9
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
2 +V
167 401 104 0 1 3
0 11
0
0 0 53488 0
2 5V
-7 -22 7 -14
3 V10
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3874 0 0
0
0
7 Pulser~
4 172 215 0 10 12
0 14 15 8 16 0 0 10 10 11
7
0
0 0 4144 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6671 0 0
0
0
5 SCOPE
12 461 66 0 1 11
0 6
0
0 0 57584 0
1 Z
-5 -4 2 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3789 0 0
0
0
5 SCOPE
12 321 66 0 1 11
0 7
0
0 0 57584 0
1 Y
-5 -4 2 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4871 0 0
0
0
5 SCOPE
12 201 66 0 1 11
0 4
0
0 0 57584 0
1 X
-5 -4 2 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3750 0 0
0
0
5 SCOPE
12 391 215 0 1 11
0 5
0
0 0 57584 0
1 W
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8778 0 0
0
0
28
0 1 5 0 0 4096 0 0 22 8 0 3
361 230
391 230
391 227
1 3 3 0 0 0 0 3 8 0 0 2
303 239
303 239
1 2 2 0 0 4224 0 4 8 0 0 4
303 230
304 230
304 230
303 230
1 1 4 0 0 0 0 6 8 0 0 2
303 221
303 221
1 5 3 0 0 4224 0 2 14 0 0 2
430 160
431 160
1 5 2 0 0 0 0 1 13 0 0 2
318 160
318 160
1 0 4 0 0 4096 0 5 0 0 15 2
206 142
201 142
0 4 5 0 0 4224 0 0 8 16 0 3
361 160
361 230
354 230
1 0 6 0 0 4112 0 9 0 0 13 2
484 78
461 78
1 0 7 0 0 4096 0 10 0 0 14 2
344 78
321 78
1 0 4 0 0 4096 0 11 0 0 15 2
224 78
201 78
1 0 8 0 0 4096 0 7 0 0 25 2
216 205
216 206
1 0 6 0 0 12288 0 19 0 0 24 4
461 78
461 77
461 77
461 142
1 0 7 0 0 0 0 20 0 0 26 2
321 78
321 85
1 6 4 0 0 4224 0 21 12 0 0 3
201 78
201 142
202 142
1 3 5 0 0 0 0 14 14 0 0 4
377 142
361 142
361 160
377 160
1 0 9 0 0 4096 0 13 0 0 18 2
264 142
249 142
0 3 9 0 0 4224 0 0 13 22 0 3
249 115
249 160
264 160
1 0 10 0 0 4096 0 12 0 0 20 2
154 142
140 142
0 3 10 0 0 4224 0 0 12 23 0 3
140 115
140 160
154 160
1 4 11 0 0 4224 0 17 14 0 0 2
401 113
401 115
1 4 9 0 0 0 0 16 13 0 0 3
249 113
249 115
288 115
1 4 10 0 0 0 0 15 12 0 0 3
140 113
140 115
178 115
6 2 6 0 0 12416 0 14 13 0 0 6
425 142
461 142
461 187
239 187
239 151
257 151
2 3 8 0 0 12416 0 14 18 0 0 4
370 151
350 151
350 206
196 206
6 2 7 0 0 12416 0 13 12 0 0 6
312 142
321 142
321 85
116 85
116 151
147 151
0 6 6 0 0 0 0 0 14 24 0 2
425 142
425 142
0 0 12 0 0 4224 0 0 0 0 0 5
297 269
568 269
568 302
297 302
297 269
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
299 266 565 303
303 270 562 298
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 25
36 265 244 289
40 269 240 285
25 Limited sequence counter.
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
