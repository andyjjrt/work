CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 432 635 647
27262994 0
0
6 Title:
5 Name:
0
0
0
53
9 Terminal~
194 17 126 0 1 3
0 2
0
0 0 49504 90
2 CN
-6 2 8 10
3 T30
-10 -25 11 -17
0
3 CN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8953 0 0
0
0
9 Terminal~
194 17 108 0 1 3
0 3
0
0 0 49504 90
1 C
-1 -14 6 -6
3 T29
-11 -25 10 -17
0
2 C;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4441 0 0
0
0
9 Terminal~
194 108 126 0 1 3
0 4
0
0 0 49504 90
2 BN
-5 3 9 11
3 T28
-10 -25 11 -17
0
3 BN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3618 0 0
0
0
9 Terminal~
194 108 108 0 1 3
0 5
0
0 0 49504 90
1 B
-1 -14 6 -6
3 T27
-11 -25 10 -17
0
2 B;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6153 0 0
0
0
9 Terminal~
194 196 126 0 1 3
0 6
0
0 0 49504 90
2 AN
-5 3 9 11
3 T26
-10 -25 11 -17
0
3 AN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5394 0 0
0
0
9 Terminal~
194 196 108 0 1 3
0 7
0
0 0 49504 90
1 A
-1 -14 6 -6
3 T25
-11 -25 10 -17
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7734 0 0
0
0
9 3-In AND~
219 505 188 0 4 22
0 7 5 3 8
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 5 0
1 U
9914 0 0
0
0
9 3-In AND~
219 505 150 0 4 22
0 6 5 3 9
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 5 0
1 U
3747 0 0
0
0
9 3-In AND~
219 505 112 0 4 22
0 7 4 3 10
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 4 0
1 U
3549 0 0
0
0
9 3-In AND~
219 505 74 0 4 22
0 6 4 3 11
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 4 0
1 U
7931 0 0
0
0
9 Terminal~
194 463 67 0 1 3
0 6
0
0 0 49504 90
2 AN
-16 -7 -2 1
3 T24
-10 -25 11 -17
0
3 AN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9325 0 0
0
0
9 Terminal~
194 463 76 0 1 3
0 4
0
0 0 49504 90
2 BN
-16 -6 -2 2
3 T23
-10 -25 11 -17
0
3 BN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8903 0 0
0
0
9 Terminal~
194 463 85 0 1 3
0 3
0
0 0 49504 90
1 C
-10 -6 -3 2
3 T22
-10 -25 11 -17
0
2 C;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3834 0 0
0
0
9 Terminal~
194 463 105 0 1 3
0 7
0
0 0 49504 90
1 A
-10 -7 -3 1
3 T21
-10 -25 11 -17
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3363 0 0
0
0
9 Terminal~
194 463 114 0 1 3
0 4
0
0 0 49504 90
2 BN
-16 -6 -2 2
3 T20
-10 -25 11 -17
0
3 BN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7668 0 0
0
0
9 Terminal~
194 463 123 0 1 3
0 3
0
0 0 49504 90
1 C
-10 -6 -3 2
3 T19
-10 -25 11 -17
0
2 C;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4718 0 0
0
0
9 Terminal~
194 463 199 0 1 3
0 3
0
0 0 49504 90
1 C
-10 -6 -3 2
3 T18
-10 -25 11 -17
0
2 C;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3874 0 0
0
0
9 Terminal~
194 463 190 0 1 3
0 5
0
0 0 49504 90
1 B
-10 -6 -3 2
3 T17
-10 -25 11 -17
0
2 B;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6671 0 0
0
0
9 Terminal~
194 463 181 0 1 3
0 7
0
0 0 49504 90
1 A
-10 -7 -3 1
3 T16
-10 -25 11 -17
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3789 0 0
0
0
9 Terminal~
194 463 161 0 1 3
0 3
0
0 0 49504 90
1 C
-10 -6 -3 2
3 T15
-10 -25 11 -17
0
2 C;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4871 0 0
0
0
9 Terminal~
194 463 152 0 1 3
0 5
0
0 0 49504 90
1 B
-10 -6 -3 2
3 T14
-10 -25 11 -17
0
2 B;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3750 0 0
0
0
9 Terminal~
194 463 143 0 1 3
0 6
0
0 0 49504 90
2 AN
-16 -7 -2 1
3 T13
-10 -25 11 -17
0
3 AN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8778 0 0
0
0
5 SCOPE
12 401 62 0 1 11
0 19
0
0 0 57568 0
3 000
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
538 0 0
0
0
5 SCOPE
12 401 100 0 1 11
0 18
0
0 0 57568 0
3 001
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6843 0 0
0
0
5 SCOPE
12 401 138 0 1 11
0 17
0
0 0 57568 0
3 010
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3136 0 0
0
0
5 SCOPE
12 401 176 0 1 11
0 16
0
0 0 57568 0
3 011
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5950 0 0
0
0
5 SCOPE
12 537 62 0 1 11
0 11
0
0 0 57568 0
3 100
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5670 0 0
0
0
5 SCOPE
12 537 100 0 1 11
0 10
0
0 0 57568 0
3 101
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6828 0 0
0
0
5 SCOPE
12 537 138 0 1 11
0 9
0
0 0 57568 0
3 110
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6735 0 0
0
0
5 SCOPE
12 537 176 0 1 11
0 8
0
0 0 57568 0
3 111
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8365 0 0
0
0
2 +V
167 94 65 0 1 3
0 13
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4132 0 0
0
0
2 +V
167 183 65 0 1 3
0 14
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4551 0 0
0
0
2 +V
167 274 65 0 1 3
0 15
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3635 0 0
0
0
7 Pulser~
4 58 165 0 10 12
0 21 22 12 23 0 0 20 20 13
8
0
0 0 4128 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3973 0 0
0
0
6 74113~
219 238 123 0 6 22
0 15 12 15 15 6 7
0
0 0 4192 512
7 74LS113
-25 -42 24 -34
3 U1A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 1 1 0
1 U
3851 0 0
0
0
6 74113~
219 149 123 0 6 22
0 14 7 14 14 4 5
0
0 0 4192 512
7 74LS113
-25 -42 24 -34
3 U1B
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 2 1 0
1 U
8383 0 0
0
0
6 74113~
219 60 123 0 6 22
0 13 5 13 13 2 3
0
0 0 4192 512
7 74LS113
-25 -42 24 -34
3 U2A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 1 2 0
1 U
9334 0 0
0
0
9 Terminal~
194 327 143 0 1 3
0 6
0
0 0 49504 90
2 AN
-16 -7 -2 1
3 T12
-10 -25 11 -17
0
3 AN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7471 0 0
0
0
9 Terminal~
194 327 152 0 1 3
0 5
0
0 0 49504 90
1 B
-10 -6 -3 2
3 T11
-10 -25 11 -17
0
2 B;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3334 0 0
0
0
9 Terminal~
194 327 161 0 1 3
0 2
0
0 0 49504 90
2 CN
-16 -6 -2 2
3 T10
-10 -25 11 -17
0
3 CN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3559 0 0
0
0
9 Terminal~
194 327 181 0 1 3
0 7
0
0 0 49504 90
1 A
-10 -7 -3 1
2 T9
-7 -25 7 -17
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
984 0 0
0
0
9 Terminal~
194 327 190 0 1 3
0 5
0
0 0 49504 90
1 B
-10 -6 -3 2
2 T8
-7 -25 7 -17
0
2 B;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7557 0 0
0
0
9 Terminal~
194 327 199 0 1 3
0 2
0
0 0 49504 90
2 CN
-16 -6 -2 2
2 T7
-7 -25 7 -17
0
3 CN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3146 0 0
0
0
9 Terminal~
194 327 123 0 1 3
0 2
0
0 0 49504 90
2 CN
-16 -6 -2 2
2 T6
-7 -25 7 -17
0
3 CN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5687 0 0
0
0
9 Terminal~
194 327 114 0 1 3
0 4
0
0 0 49504 90
2 BN
-16 -6 -2 2
2 T5
-7 -25 7 -17
0
3 BN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
7939 0 0
0
0
9 Terminal~
194 327 105 0 1 3
0 7
0
0 0 49504 90
1 A
-10 -7 -3 1
2 T4
-7 -25 7 -17
0
2 A;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3308 0 0
0
0
9 Terminal~
194 327 85 0 1 3
0 2
0
0 0 49504 90
2 CN
-16 -6 -2 2
2 T3
-7 -25 7 -17
0
3 CN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3408 0 0
0
0
9 Terminal~
194 327 76 0 1 3
0 4
0
0 0 49504 90
2 BN
-16 -6 -2 2
2 T2
-7 -25 7 -17
0
3 BN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
9773 0 0
0
0
9 Terminal~
194 327 67 0 1 3
0 6
0
0 0 49504 90
2 AN
-16 -7 -2 1
2 T1
-7 -25 7 -17
0
3 AN;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
691 0 0
0
0
9 3-In AND~
219 369 74 0 4 22
0 6 4 2 19
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 3 0
1 U
7834 0 0
0
0
9 3-In AND~
219 369 112 0 4 22
0 7 4 2 18
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 3 0
1 U
3588 0 0
0
0
9 3-In AND~
219 369 150 0 4 22
0 6 5 2 17
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U3C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 3 0
1 U
4528 0 0
0
0
9 3-In AND~
219 369 188 0 4 22
0 7 5 2 16
0
0 0 96 0
6 74LS11
-21 -28 21 -20
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 4 0
1 U
3303 0 0
0
0
51
0 0 20 0 0 16 0 0 0 0 0 5
305 264
576 264
576 296
305 296
305 264
1 5 2 0 0 0 0 1 37 0 0 2
28 124
28 124
1 6 3 0 0 4096 0 2 37 0 0 2
28 106
34 106
1 5 4 0 0 4096 0 3 36 0 0 2
119 124
117 124
1 0 5 0 0 0 0 4 0 0 24 2
119 106
119 106
1 5 6 0 0 4096 0 5 35 0 0 2
207 124
206 124
1 0 7 0 0 0 0 6 0 0 25 2
207 106
207 106
1 4 8 0 0 4224 0 30 7 0 0 2
537 188
526 188
1 4 9 0 0 4224 0 29 8 0 0 2
537 150
526 150
1 4 10 0 0 4224 0 28 9 0 0 2
537 112
526 112
1 4 11 0 0 4224 0 27 10 0 0 2
537 74
526 74
1 3 3 0 0 4224 0 17 7 0 0 2
474 197
481 197
1 2 5 0 0 4096 0 18 7 0 0 2
474 188
481 188
1 1 7 0 0 4096 0 19 7 0 0 2
474 179
481 179
1 3 3 0 0 0 0 20 8 0 0 2
474 159
481 159
1 2 5 0 0 0 0 21 8 0 0 2
474 150
481 150
1 1 6 0 0 4224 0 22 8 0 0 2
474 141
481 141
1 3 3 0 0 0 0 16 9 0 0 2
474 121
481 121
1 2 4 0 0 4224 0 15 9 0 0 2
474 112
481 112
1 1 7 0 0 4096 0 14 9 0 0 4
474 103
482 103
482 103
481 103
1 3 3 0 0 0 0 13 10 0 0 2
474 83
481 83
1 2 4 0 0 0 0 12 10 0 0 2
474 74
481 74
1 1 6 0 0 0 0 11 10 0 0 2
474 65
481 65
2 6 5 0 0 4224 0 37 36 0 0 4
89 115
119 115
119 106
123 106
2 6 7 0 0 4224 0 36 35 0 0 4
178 115
207 115
207 106
212 106
2 3 12 0 0 8320 0 35 34 0 0 3
267 115
267 156
82 156
1 0 13 0 0 4096 0 37 0 0 29 2
82 106
94 106
4 0 13 0 0 4096 0 37 0 0 29 2
58 79
94 79
3 1 13 0 0 8320 0 37 31 0 0 3
82 124
94 124
94 74
4 0 14 0 0 4096 0 36 0 0 32 2
147 79
183 79
1 0 14 0 0 0 0 36 0 0 32 2
171 106
183 106
1 3 14 0 0 4224 0 32 36 0 0 3
183 74
183 124
171 124
4 0 15 0 0 4096 0 35 0 0 35 2
236 79
274 79
1 0 15 0 0 0 0 35 0 0 35 2
260 106
274 106
1 3 15 0 0 4224 0 33 35 0 0 3
274 74
274 124
260 124
1 4 16 0 0 4224 0 26 53 0 0 2
401 188
390 188
1 4 17 0 0 4224 0 25 52 0 0 2
401 150
390 150
1 4 18 0 0 4224 0 24 51 0 0 2
401 112
390 112
1 4 19 0 0 4224 0 23 50 0 0 2
401 74
390 74
1 3 2 0 0 4224 0 43 53 0 0 2
338 197
345 197
1 2 5 0 0 0 0 42 53 0 0 2
338 188
345 188
1 1 7 0 0 0 0 41 53 0 0 2
338 179
345 179
1 3 2 0 0 0 0 40 52 0 0 2
338 159
345 159
1 2 5 0 0 0 0 39 52 0 0 2
338 150
345 150
1 1 6 0 0 0 0 38 52 0 0 2
338 141
345 141
1 3 2 0 0 0 0 44 51 0 0 2
338 121
345 121
1 2 4 0 0 0 0 45 51 0 0 2
338 112
345 112
1 1 7 0 0 0 0 46 51 0 0 4
338 103
346 103
346 103
345 103
1 3 2 0 0 0 0 47 50 0 0 2
338 83
345 83
1 2 4 0 0 0 0 48 50 0 0 2
338 74
345 74
1 1 6 0 0 0 0 49 50 0 0 2
338 65
345 65
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
307 261 573 298
311 265 570 293
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 45
24 258 256 302
28 262 252 294
45 Using AND gates to decode a 
MOD-8 counter.
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
