CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 390
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 390 635 516
25165842 0
0
6 Title:
5 Name:
0
0
0
10
5 SCOPE
12 162 15 0 1 11
0 12
0
0 0 57568 0
1 D
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SCOPE
12 200 15 0 1 11
0 11
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 491 19 0 1 11
0 9
0
0 0 57568 0
2 QD
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 350 18 0 1 11
0 10
0
0 0 57568 0
3 QJK
-11 -4 10 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
7 Ground~
168 319 146 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 288 79 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
5 4027~
219 319 132 0 7 32
0 2 12 11 13 2 14 10
0
0 0 4192 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 512 2 1 1 0
1 U
9914 0 0
0
0
9 Inverter~
13 251 114 0 2 22
0 12 13
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3747 0 0
0
0
9 Data Seq~
170 103 43 0 17 18
0 15 16 17 18 19 20 12 11 21
22 1 1 32 5 6 0 33
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
3549 0 0
0
0
AAAAABACADAAABACADAAABACADAAABACADAAABACADAAABACADAAABACADAAABACAD
12 D Flip-Flop~
219 459 113 0 4 9
0 12 11 23 9
0
0 0 4192 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
18
0 0 3 0 0 16 0 0 0 0 0 5
309 220
580 220
580 252
309 252
309 220
0 0 4 0 0 4224 0 0 0 0 0 2
375 81
394 81
0 0 5 0 0 4224 0 0 0 0 0 2
375 91
394 91
0 0 6 0 0 4224 0 0 0 0 0 2
375 86
394 86
0 0 7 0 0 12672 0 0 0 0 0 5
408 55
503 55
503 117
406 117
406 55
0 0 8 0 0 4480 0 0 0 0 0 5
223 56
362 56
362 160
223 160
223 56
1 4 9 0 0 4224 0 3 10 0 0 3
491 31
491 77
483 77
1 7 10 0 0 4224 0 4 7 0 0 3
350 30
350 96
343 96
1 0 11 0 0 4096 0 2 0 0 17 2
200 27
200 45
1 0 12 0 0 4096 0 1 0 0 15 2
162 27
162 36
1 1 2 0 0 8320 0 6 7 0 0 4
288 73
288 68
319 68
319 75
1 5 2 0 0 0 0 5 7 0 0 2
319 140
319 138
2 0 12 0 0 4096 0 7 0 0 14 2
295 96
234 96
1 0 12 0 0 8192 0 8 0 0 15 3
236 114
234 114
234 36
7 1 12 0 0 12416 0 9 10 0 0 6
135 70
162 70
162 36
427 36
427 77
435 77
0 2 11 0 0 4224 0 0 10 17 0 4
271 45
418 45
418 95
435 95
3 8 11 0 0 0 0 7 9 0 0 6
295 105
271 105
271 45
200 45
200 79
135 79
2 4 13 0 0 4224 0 8 7 0 0 2
272 114
295 114
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 69
24 209 248 273
28 213 244 261
69 Edge-triggered D flip-flop 
implementation from a J-K 
flip-flop.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
311 217 577 254
315 221 574 249
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
276 161 308 185
280 165 304 181
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
443 161 475 185
447 165 471 181
3 (b)
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
