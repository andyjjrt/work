CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 396
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 396 635 522
27262994 0
0
6 Title:
5 Name:
0
0
0
7
5 SCOPE
12 245 118 0 1 11
0 6
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SCOPE
12 280 118 0 1 11
0 5
0
0 0 57568 0
1 S
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 315 118 0 1 11
0 4
0
0 0 57568 0
1 R
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 458 95 0 1 11
0 3
0
0 0 57568 0
1 Q
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
9 Data Seq~
170 186 122 0 17 18
0 8 9 10 11 12 4 5 6 13
14 11 1 100 2 2 0 101
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
5394 0 0
0
0
AAAEAGAGAGAGAHAHAHAHAHAGAGAEAEAGAHAHAHAHAHAGAGAGAGAGAHAHAHAHAHAGAGAGAGACADADADAD
ADACAGAGAGAGAHAHAHAHAHAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAG
AGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAGAG
6 74112~
219 413 159 0 7 32
0 5 7 6 7 4 15 3
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 1 0
1 U
7734 0 0
0
0
2 +V
167 376 108 0 1 3
0 7
0
0 0 53600 0
3 +5V
-10 -13 11 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
10
0 0 2 0 0 16 0 0 0 0 0 5
328 228
599 228
599 261
328 261
328 228
1 7 3 0 0 8320 0 4 6 0 0 3
458 107
458 123
437 123
1 0 4 0 0 4096 0 3 0 0 6 2
315 130
315 140
1 0 5 0 0 4096 0 2 0 0 7 2
280 130
280 149
1 0 6 0 0 4096 0 1 0 0 8 2
245 130
245 158
5 6 4 0 0 16512 0 6 5 0 0 5
413 171
413 175
348 175
348 140
218 140
1 7 5 0 0 16512 0 6 5 0 0 5
413 96
413 90
357 90
357 149
218 149
3 8 6 0 0 12416 0 6 5 0 0 4
383 132
366 132
366 158
218 158
2 0 7 0 0 4096 0 6 0 0 10 2
389 123
376 123
4 1 7 0 0 8320 0 6 7 0 0 3
389 141
376 141
376 117
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 80
11 217 307 281
15 221 303 269
80 Waveforms showing how a clocked 
flip-flop responds to asynchronous 
inputs.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
330 225 596 262
334 229 593 257
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 2
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
