CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 541
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 541
8388626 0
0
6 Title:
5 Name:
0
0
0
18
5 4049~
219 181 299 0 2 22
0 7 6
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U2D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 4 2 0
1 U
8953 0 0
0
0
5 4081~
219 344 317 0 3 22
0 4 3 2
0
0 0 96 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 5 0
1 U
4441 0 0
0
0
14 Logic Display~
6 391 279 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
5 4071~
219 232 308 0 3 22
0 6 5 4
0
0 0 96 0
4 4071
-7 -24 21 -16
3 U6A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 6 0
1 U
6153 0 0
0
0
13 Logic Switch~
5 299 326 0 1 11
0 3
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
1 A
-23 -3 -16 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 134 317 0 1 11
0 5
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
1 C
-23 -3 -16 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 134 299 0 1 11
0 7
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
1 B
-23 -3 -16 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 78 125 0 1 11
0 9
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 C
-24 -3 -17 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 78 221 0 1 11
0 10
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 B
-24 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 78 89 0 1 11
0 8
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-24 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7931 0 0
0
0
5 4073~
219 241 212 0 4 22
0 8 9 10 14
0
0 0 96 0
4 4073
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
9325 0 0
0
0
5 4049~
219 177 89 0 2 22
0 8 12
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 2 2 0
1 U
8903 0 0
0
0
5 4049~
219 258 156 0 2 22
0 10 15
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 2 0
1 U
3834 0 0
0
0
5 4049~
219 177 125 0 2 22
0 9 11
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U2C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 3 2 0
1 U
3363 0 0
0
0
14 Logic Display~
6 460 96 0 1 2
10 17
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7668 0 0
0
0
5 4073~
219 317 116 0 4 22
0 13 8 15 16
0
0 0 96 0
4 4073
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 4 0
1 U
4718 0 0
0
0
5 4071~
219 398 125 0 3 22
0 16 14 17
0
0 0 96 0
4 4071
-7 -24 21 -16
3 U6B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 6 0
1 U
3874 0 0
0
0
5 4011~
219 241 107 0 3 22
0 12 11 13
0
0 0 96 0
4 4011
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 3 0
1 U
6671 0 0
0
0
20
1 3 2 0 0 16 0 3 2 0 0 3
391 297
391 317
365 317
2 1 3 0 0 16 0 2 5 0 0 2
320 326
311 326
1 3 4 0 0 16 0 2 4 0 0 2
320 308
265 308
2 1 5 0 0 16 0 4 6 0 0 2
219 317
146 317
1 2 6 0 0 16 0 4 1 0 0 2
219 299
202 299
1 1 7 0 0 16 0 1 7 0 0 2
166 299
146 299
2 0 8 0 0 12416 0 16 0 0 8 5
293 116
284 116
284 66
142 66
142 89
1 0 8 0 0 0 0 11 0 0 11 3
217 203
142 203
142 89
2 0 9 0 0 4224 0 11 0 0 15 3
217 212
124 212
124 125
1 0 10 0 0 8192 0 13 0 0 16 3
243 156
191 156
191 221
1 1 8 0 0 0 0 12 10 0 0 2
162 89
90 89
2 2 11 0 0 12416 0 18 14 0 0 4
217 116
209 116
209 125
198 125
1 2 12 0 0 12416 0 18 12 0 0 4
217 98
208 98
208 89
198 89
1 3 13 0 0 4224 0 16 18 0 0 2
293 107
268 107
1 1 9 0 0 0 0 14 8 0 0 2
162 125
90 125
3 1 10 0 0 4224 0 11 9 0 0 2
217 221
90 221
2 4 14 0 0 12416 0 17 11 0 0 4
385 134
360 134
360 212
262 212
3 2 15 0 0 8320 0 16 13 0 0 4
293 125
284 125
284 156
279 156
1 4 16 0 0 4224 0 17 16 0 0 2
385 116
338 116
1 3 17 0 0 8320 0 15 17 0 0 3
460 114
460 125
431 125
25
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 124
34 384 554 428
38 388 550 420
124 Algebraic Simplification. It is obvious that the circuit in (b) 
is a great deal simpler than the original circuit in (a).
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
264 286 296 310
268 290 292 306
3 B+C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
356 319 428 343
360 323 424 339
8 z=A(B+C)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
255 347 287 371
259 351 283 367
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
388 311 404 335
392 315 400 331
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
253 231 285 255
257 235 281 251
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
262 45 286 69
266 49 282 65
2 AC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
267 160 283 184
271 164 279 180
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
269 106 285 130
273 110 281 126
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
267 145 283 169
271 149 279 165
1 _
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
262 26 286 50
266 30 282 46
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
417 131 521 155
421 135 517 151
12 z=ABC+AB(AC)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
331 93 387 117
335 97 383 113
6 AB(AC)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
206 184 222 208
210 188 218 204
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
498 123 514 147
502 127 510 143
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
489 123 505 147
493 127 501 143
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
489 113 513 137
493 117 509 133
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
364 84 380 108
368 88 376 104
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
355 84 371 108
359 88 367 104
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
356 74 380 98
360 78 376 94
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
473 123 489 147
477 127 485 143
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
339 85 355 109
343 89 351 105
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
262 36 278 60
266 40 274 56
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
270 36 286 60
274 40 282 56
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
259 193 291 217
263 197 287 213
3 ABC
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
