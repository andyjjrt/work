CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
2 70 633 528
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
2 70 633 528
8912914 0
0
6 Title:
5 Name:
0
0
0
14
13 Logic Switch~
5 125 92 0 1 11
0 16
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
6 MSB  D
-59 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 125 127 0 1 11
0 15
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
1 C
-24 -5 -17 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 125 159 0 1 11
0 14
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
1 B
-23 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 126 193 0 1 11
0 13
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
6 LSB  A
-59 -3 -17 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
9 Terminal~
194 298 148 0 1 3
0 2
0
0 0 49504 270
4 VOUT
4 -5 32 3
2 T1
-7 -25 7 -17
0
5 VOUT;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5394 0 0
0
0
7 Ground~
168 202 207 0 1 3
0 3
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
2 +V
167 236 175 0 1 3
0 17
0
0 0 54368 180
4 -15V
0 -2 28 6
2 V2
7 -12 21 -4
3 -Vs
-10 -1 11 7
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
2 +V
167 236 126 0 1 3
0 18
0
0 0 54368 0
3 15V
-10 -22 11 -14
2 V1
-7 -32 7 -24
3 +Vs
-11 -14 10 -6
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
8 Op-Amp5~
219 236 147 0 5 11
0 3 12 18 17 2
0
0 0 1088 0
6 OPAMP5
16 -25 58 -17
2 U1
30 -35 44 -27
6 Op amp
5 9 47 17
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
9 Resistor~
219 155 92 0 2 5
0 16 12
0
0 0 352 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 155 127 0 2 5
0 15 12
0
0 0 352 0
2 2k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 154 159 0 2 5
0 14 12
0
0 0 352 0
2 4k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 155 193 0 2 5
0 13 12
0
0 0 352 0
2 8k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 233 92 0 2 5
0 12 2
0
0 0 864 0
2 1k
-7 -14 7 -6
2 Rf
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
23
0 0 4 0 0 8320 0 0 0 0 0 8
375 32
375 28
408 28
408 23
408 23
408 28
439 28
439 32
0 0 5 0 0 24704 0 0 0 0 0 8
65 208
65 214
100 214
100 221
100 221
100 214
137 214
137 208
0 0 6 0 0 4224 0 0 0 0 0 2
370 36
546 36
0 0 7 0 0 4224 0 0 0 0 0 2
370 307
546 307
0 0 8 0 0 4224 0 0 0 0 0 2
370 244
546 244
0 0 9 0 0 4224 0 0 0 0 0 2
370 180
546 180
0 0 10 0 0 4224 0 0 0 0 0 2
370 115
546 115
0 0 11 0 0 4224 0 0 0 0 0 2
370 52
546 52
0 0 1 0 0 4256 0 0 0 0 0 2
447 39
447 304
2 0 2 0 0 8320 0 14 0 0 11 3
251 92
268 92
268 147
5 1 2 0 0 0 0 9 5 0 0 2
254 147
286 147
1 0 12 0 0 8192 0 14 0 0 14 3
215 92
202 92
202 141
1 1 3 0 0 8320 0 9 6 0 0 3
218 153
202 153
202 201
2 0 12 0 0 0 0 9 0 0 17 2
218 141
181 141
2 0 12 0 0 0 0 11 0 0 17 2
173 127
181 127
2 0 12 0 0 0 0 12 0 0 17 2
172 159
181 159
2 2 12 0 0 8320 0 10 13 0 0 4
173 92
181 92
181 193
173 193
1 1 13 0 0 4224 0 4 13 0 0 2
138 193
137 193
1 1 14 0 0 4224 0 3 12 0 0 2
137 159
136 159
1 1 15 0 0 0 0 2 11 0 0 2
137 127
137 127
1 1 16 0 0 0 0 1 10 0 0 2
137 92
137 92
1 4 17 0 0 0 0 7 9 0 0 2
236 160
236 160
1 3 18 0 0 4224 0 8 9 0 0 2
236 135
236 134
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 79
102 360 470 404
106 364 466 396
79 Simple DAC using an op-amp summing amplifier 
with binary-weighted resistors.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 170
451 31 555 375
455 35 551 307
170 VOUT (volts)
     0
  -0.625
  -1.250
  -1.875
  -2.500
  -3.125
  -3.750
  -4.375
  -5.000
  -5.625
  -6.250
  -6.875
  -7.500
  -8.125
  -8.750
  -9.375
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 49
427 32 451 376
431 36 447 308
49 A
0
1
0
1
0
1
0
1
0
1
0
1
0
1
0
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 49
409 32 433 376
413 36 429 308
49 B
0
0
1
1
0
0
1
1
0
0
1
1
0
0
1
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 49
390 32 414 376
394 36 410 308
49 C
0
0
0
0
1
1
1
1
0
0
0
0
1
1
1
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 49
371 32 395 376
375 36 391 308
49 D
0
0
0
0
0
0
0
0
1
1
1
1
1
1
1
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
524 63 556 87
528 67 552 83
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
524 287 556 311
528 291 552 307
3 MSB
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
370 3 447 23
374 7 444 21
10 Input Code
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 25
47 222 159 259
51 226 156 254
25 Digital inputs:
0V or 5V
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
440 319 472 343
444 323 468 339
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
177 319 209 343
181 323 205 339
3 (a)
0
1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
438174074 1210432 100 100 0 0
77 66 587 216
7 94 168 164
587 66
77 66
587 66
587 216
0 0
0.01 0 0.01 1.05685e-314 0.01 0.01
12401 0
4 1 10
1
280 147
0 2 0 0 1	0 11 0 0
829752294 8550464 100 100 0 0
77 66 587 246
4 405 625 740
586 66
77 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 1e-006 10
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
