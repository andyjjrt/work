CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 436 635 561
27262994 0
0
6 Title:
5 Name:
0
0
0
16
7 Ground~
168 82 126 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8953 0 0
0
0
12 Hex Display~
7 91 72 0 16 19
10 5 4 3 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4441 0 0
0
0
6 74113~
219 191 179 0 6 22
0 9 6 9 9 13 3
0
0 0 4192 512
7 74LS113
-25 -42 24 -34
3 U2A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 2 0
1 U
3618 0 0
0
0
6 74113~
219 280 179 0 6 22
0 10 7 10 10 6 4
0
0 0 4192 512
7 74LS113
-25 -42 24 -34
3 U1B
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 2 1 0
1 U
6153 0 0
0
0
6 74113~
219 369 179 0 6 22
0 11 8 11 11 7 5
0
0 0 4192 512
7 74LS113
-25 -42 24 -34
3 U1A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 1 1 0
1 U
5394 0 0
0
0
14 Logic Display~
6 357 74 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 268 74 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 176 74 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
7 Pulser~
4 464 180 0 10 12
0 14 15 8 16 0 0 20 20 21
7
0
0 0 4128 512
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3549 0 0
0
0
5 SCOPE
12 428 80 0 1 11
0 8
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
5 SCOPE
12 334 80 0 1 11
0 5
0
0 0 57568 0
1 A
-4 -4 3 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
5 SCOPE
12 245 80 0 1 11
0 4
0
0 0 57568 0
1 B
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
5 SCOPE
12 153 80 0 1 11
0 3
0
0 0 57568 0
1 C
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
2 +V
167 405 121 0 1 3
0 11
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
2 +V
167 314 121 0 1 3
0 10
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
2 +V
167 225 121 0 1 3
0 9
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
24
0 0 12 0 0 16 0 0 0 0 0 5
306 272
577 272
577 304
306 304
306 272
4 1 2 0 0 4224 0 2 1 0 0 2
82 96
82 120
3 0 3 0 0 8192 0 2 0 0 11 3
88 96
88 113
153 113
2 0 4 0 0 8320 0 2 0 0 12 3
94 96
94 107
245 107
1 0 5 0 0 8320 0 2 0 0 13 3
100 96
100 101
334 101
2 5 6 0 0 4224 0 3 4 0 0 4
220 171
235 171
235 180
248 180
2 5 7 0 0 4224 0 4 5 0 0 4
309 171
325 171
325 180
337 180
1 0 3 0 0 0 0 8 0 0 11 2
176 92
153 92
1 0 4 0 0 0 0 7 0 0 12 2
268 92
245 92
1 0 5 0 0 0 0 6 0 0 13 2
357 92
334 92
1 6 3 0 0 4224 0 13 3 0 0 3
153 92
153 162
165 162
1 6 4 0 0 0 0 12 4 0 0 3
245 92
245 162
254 162
1 6 5 0 0 0 0 11 5 0 0 3
334 92
334 162
343 162
1 0 8 0 0 4224 0 10 0 0 15 2
428 92
428 171
3 2 8 0 0 0 0 9 5 0 0 2
440 171
398 171
1 0 9 0 0 4096 0 3 0 0 18 2
213 162
225 162
4 0 9 0 0 4096 0 3 0 0 18 2
189 135
225 135
3 1 9 0 0 8320 0 3 16 0 0 3
213 180
225 180
225 130
4 0 10 0 0 4096 0 4 0 0 21 2
278 135
314 135
1 0 10 0 0 0 0 4 0 0 21 2
302 162
314 162
1 3 10 0 0 4224 0 15 4 0 0 3
314 130
314 180
302 180
4 0 11 0 0 4096 0 5 0 0 24 2
367 135
405 135
1 0 11 0 0 0 0 5 0 0 24 2
391 162
405 162
1 3 11 0 0 4224 0 14 5 0 0 3
405 130
405 180
391 180
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
308 269 574 306
312 273 571 301
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 19
42 279 202 303
46 283 198 299
19 MOD-8 down counter.
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
