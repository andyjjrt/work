CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 485
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 485 635 577
25165842 0
0
6 Title:
5 Name:
0
0
0
11
5 SCOPE
12 529 169 0 1 11
0 4
0
0 0 57584 0
2 CP
-8 -4 6 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
7 Pulser~
4 463 245 0 10 12
0 18 19 4 20 0 0 5 5 6
7
0
0 0 1072 0
0
2 V2
-7 -28 7 -20
5 Clock
-17 20 18 28
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 1 0 0
1 V
4441 0 0
0
0
2 +V
167 499 134 0 1 3
0 7
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
6 74113~
219 464 193 0 6 22
0 7 4 7 7 21 6
0
0 0 4208 512
7 74LS113
-25 -42 24 -34
3 U3A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 1 0
1 U
6153 0 0
0
0
6 74113~
219 381 193 0 6 22
0 7 6 7 7 22 5
0
0 0 4208 512
7 74LS113
-25 -42 24 -34
3 U3B
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 2 1 0
1 U
5394 0 0
0
0
6 74113~
219 296 193 0 6 22
0 7 5 7 7 23 9
0
0 0 4208 512
7 74LS113
-25 -42 24 -34
3 U4A
-13 24 8 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 2 0
1 U
7734 0 0
0
0
5 SCOPE
12 258 55 0 1 11
0 8
0
0 0 57584 0
1 Z
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
7 Ground~
168 243 148 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 62 160 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
6 PROM32
80 109 117 0 14 29
0 2 2 2 2 2 2 17 16 15
14 13 12 11 10
0
0 0 1392 692
7 Storage
-25 45 24 53
2 U2
-7 -61 7 -53
8 register
-28 56 28 64
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 2 3 4 5 6 7 9 10
11 12 13 14 15 1 2 3 4 5
6 7 9 10 11 12 13 14 15 0
65 0 0 0 1 1 0 0
1 U
7931 0 0
0
0
LFAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
7 74LS151
20 200 117 0 14 29
0 17 16 15 14 13 12 11 10 2
9 5 6 8 24
0
0 0 12528 692
7 74HC151
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
33
0 0 3 0 0 4224 0 0 0 0 0 5
319 307
590 307
590 340
319 340
319 307
1 0 4 0 0 4096 0 1 0 0 3 2
529 181
529 185
3 2 4 0 0 8320 0 2 4 0 0 4
487 236
529 236
529 185
493 185
2 6 5 0 0 4096 0 6 5 0 0 4
325 185
347 185
347 176
355 176
2 6 6 0 0 4096 0 5 4 0 0 4
410 185
430 185
430 176
438 176
1 0 7 0 0 4096 0 6 0 0 7 2
318 176
331 176
3 0 7 0 0 8192 0 6 0 0 12 3
318 194
331 194
331 146
1 0 7 0 0 0 0 5 0 0 9 2
403 176
416 176
3 0 7 0 0 0 0 5 0 0 12 3
403 194
416 194
416 146
4 0 7 0 0 0 0 5 0 0 12 2
379 149
379 146
4 0 7 0 0 0 0 4 0 0 12 2
462 149
462 146
4 0 7 0 0 8320 0 6 0 0 14 3
294 149
294 146
499 146
1 0 7 0 0 0 0 4 0 0 14 2
486 176
499 176
1 3 7 0 0 0 0 3 4 0 0 3
499 143
499 194
486 194
1 13 8 0 0 8320 0 7 11 0 0 3
258 67
258 82
232 82
6 10 9 0 0 8320 0 6 11 0 0 4
270 176
261 176
261 127
232 127
0 11 5 0 0 8320 0 0 11 4 0 3
347 176
347 118
232 118
0 12 6 0 0 8320 0 0 11 5 0 3
430 176
430 109
232 109
1 9 2 0 0 4096 0 8 11 0 0 3
243 142
243 136
238 136
5 0 2 0 0 4096 0 10 0 0 25 2
77 82
62 82
4 0 2 0 0 0 0 10 0 0 25 2
77 91
62 91
3 0 2 0 0 0 0 10 0 0 25 2
77 100
62 100
2 0 2 0 0 0 0 10 0 0 25 2
77 109
62 109
1 0 2 0 0 0 0 10 0 0 25 2
71 145
62 145
6 1 2 0 0 8320 0 10 9 0 0 3
77 73
62 73
62 154
14 8 10 0 0 4224 0 10 11 0 0 2
141 73
168 73
13 7 11 0 0 4224 0 10 11 0 0 2
141 82
168 82
12 6 12 0 0 4224 0 10 11 0 0 2
141 91
168 91
11 5 13 0 0 4224 0 10 11 0 0 2
141 100
168 100
10 4 14 0 0 4224 0 10 11 0 0 2
141 109
168 109
9 3 15 0 0 4224 0 10 11 0 0 2
141 118
168 118
8 2 16 0 0 4224 0 10 11 0 0 2
141 127
168 127
7 1 17 0 0 4224 0 10 11 0 0 2
141 136
168 136
5
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
172 154 228 191
176 158 225 186
14 8-input
  MUX
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
133 133 154 153
137 137 151 151
2 X7
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
133 55 154 75
137 59 151 73
2 X0
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 77
30 297 278 361
34 301 274 349
77 Parallel-to-serial converter. 
Storage register contains
X7-X0 = 10110101.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
321 304 587 341
325 308 584 336
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
267780172 8525888 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.0159882 0 5.36094e-315 0 0.016 0.016
12401 0
4 1e-006 2
2
221 112
0 7 0 0 2	0 34 0 0
367 106
0 2 0 0 1	0 34 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 34 0 0
200 112
0 7 0 0 2	0 34 0 0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
