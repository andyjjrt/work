CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 418
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 418
11010070 0
0
6 Title:
5 Name:
0
0
0
11
9 Terminal~
194 179 140 0 1 3
0 2
0
0 0 49520 90
6 OUTPUT
-50 -5 -8 3
2 T1
-7 -25 7 -17
0
7 OUTPUT;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8953 0 0
0
0
7 Ground~
168 254 232 0 1 3
0 3
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4441 0 0
0
0
7 Ground~
168 337 232 0 1 3
0 3
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 386 232 0 1 3
0 3
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
2 +V
167 386 51 0 1 3
0 5
0
0 0 53616 0
3 +5V
-11 -14 10 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
10 Capacitor~
219 337 206 0 2 5
0 7 3
0
0 0 336 270
5 .01uF
-46 -3 -11 5
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
10 Capacitor~
219 386 206 0 2 5
0 4 3
0
0 0 592 270
5 .01uF
5 8 40 16
1 C
14 -3 21 5
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
10 555 Timer~
219 295 129 0 8 17
0 3 4 2 5 7 4 6 5
0
0 0 12496 0
3 555
-11 -36 10 -28
2 U1
-7 -46 7 -38
0
0
29 %D %1 %2 %3 %4 %5 %6 %7 %8 %S
0
0
4 CAN8
17

0 1 2 3 4 5 6 7 8 1
2 3 4 5 6 7 8 0
88 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
4 .IC~
207 295 172 0 1 3
0 4
0
0 0 53328 0
2 5V
-7 -16 7 -8
4 CMD1
-14 -26 14 -18
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
3549 0 0
0
0
9 Resistor~
219 386 155 0 2 5
0 6 4
0
0 0 624 270
4 100k
1 0 29 8
2 RB
8 -5 22 3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 386 96 0 3 5
0 5 6 1
0
0 0 624 270
3 10k
5 0 26 8
2 RA
8 -5 22 3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
14
1 0 4 0 0 0 0 9 0 0 9 2
295 184
295 184
1 2 3 0 0 4096 0 4 7 0 0 2
386 226
386 215
1 2 3 0 0 0 0 3 6 0 0 2
337 226
337 215
3 1 2 0 0 4224 0 8 1 0 0 2
263 138
190 138
8 0 5 0 0 8192 0 8 0 0 6 3
327 120
336 120
336 68
4 0 5 0 0 12416 0 8 0 0 8 4
263 147
231 147
231 68
386 68
1 1 3 0 0 8320 0 8 2 0 0 3
263 120
254 120
254 226
1 1 5 0 0 0 0 5 11 0 0 2
386 60
386 78
2 0 4 0 0 12416 0 8 0 0 10 4
263 129
243 129
243 184
348 184
6 0 4 0 0 0 0 8 0 0 13 4
327 138
348 138
348 184
386 184
7 0 6 0 0 4224 0 8 0 0 14 2
327 129
386 129
5 1 7 0 0 8320 0 8 6 0 0 3
327 147
337 147
337 197
2 1 4 0 0 0 0 10 7 0 0 2
386 173
386 197
2 1 6 0 0 0 0 11 10 0 0 2
386 114
386 137
1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 46
110 267 486 291
114 271 482 287
46 555 timer IC used as an astable multivibrator.
63 .OPTIONS ITL1=1000 ITL4=100 RELTOL=0.01 CONVLIMIT RSHUNT=1E12

16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.006 1e-005 1e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
625541492 8550464 100 100 0 0
77 66 587 156
4 418 635 639
587 66
77 66
587 66
587 156
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 0.001 2
2
207 138
0 2 0 0 1	0 4 0 0
365 184
0 4 0 0 3	0 10 0 0
47318444 8550464 100 100 0 0
77 66 587 156
4 418 635 639
586 66
77 66
587 66
587 156
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 1e-006 2
2
219 152
0 3 0 0 1	0 5 0 0
378 198
0 4 0 0 3	0 11 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
