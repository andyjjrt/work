CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
2 70 633 462
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
2 70 633 462
8912914 0
0
6 Title:
5 Name:
0
0
0
34
13 Logic Switch~
5 321 275 0 1 11
0 17
0
0 0 21600 602
2 0V
11 0 25 8
2 V5
11 -10 25 -2
9 B3  (MSB)
-7 16 56 24
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 263 274 0 1 11
0 18
0
0 0 21600 602
2 0V
11 0 25 8
2 V4
11 -10 25 -2
2 B2
-6 16 8 24
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 206 275 0 1 11
0 19
0
0 0 21600 602
2 0V
11 0 25 8
2 V3
11 -10 25 -2
2 B1
-7 15 7 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 149 276 0 1 11
0 20
0
0 0 21600 602
2 0V
11 0 25 8
2 V2
11 -10 25 -2
9 (LSB)  B0
-56 15 7 23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
7 Buffer~
58 320 248 0 2 22
0 17 4
0
0 0 96 90
4 4050
-14 -19 14 -11
3 U2D
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 4 1 0
1 U
5394 0 0
0
0
7 Buffer~
58 262 248 0 2 22
0 18 5
0
0 0 96 90
4 4050
-14 -19 14 -11
3 U2C
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 3 1 0
1 U
7734 0 0
0
0
7 Buffer~
58 205 248 0 2 22
0 19 6
0
0 0 96 90
4 4050
-14 -19 14 -11
3 U2B
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 2 1 0
1 U
9914 0 0
0
0
9 Terminal~
194 477 184 0 1 3
0 2
0
0 0 49504 270
4 VOUT
4 -5 32 3
2 T1
-7 -25 7 -17
0
5 VOUT;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3747 0 0
0
0
7 Ground~
168 364 208 0 1 3
0 3
0
0 0 53344 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3549 0 0
0
0
2 +V
167 102 85 0 1 3
0 16
0
0 0 54368 90
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
5 +VREF
-41 -6 -6 2
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
7 Ground~
168 103 192 0 1 3
0 3
0
0 0 53344 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
11 Contacts:B~
215 326 110 0 10 18
0 8 16 3 0 0 0 0 0 0
1
0
0 0 96 782
6 NORMAL
-19 -25 23 -17
4 RLY5
-12 -35 16 -27
2 B3
-5 -45 9 -37
0
17 %D %1 %2 %3 %I %S
0
15 alias:XCONTACTS
4 SIP3
7

0 1 2 3 1 2 3 0
88 0 0 0 1 0 -5 0
3 RLY
8903 0 0
0
0
7 Ground~
168 356 113 0 1 3
0 3
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
11 Contacts:B~
215 269 110 0 10 18
0 9 16 3 0 0 0 0 0 0
1
0
0 0 96 782
6 NORMAL
-19 -25 23 -17
4 RLY4
-12 -35 16 -27
2 B2
-5 -45 9 -37
0
17 %D %1 %2 %3 %I %S
0
15 alias:XCONTACTS
4 SIP3
7

0 1 2 3 1 2 3 0
88 0 0 0 1 0 -4 0
3 RLY
3363 0 0
0
0
7 Ground~
168 299 113 0 1 3
0 3
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7668 0 0
0
0
11 Contacts:B~
215 212 110 0 10 18
0 10 16 3 0 0 0 0 0 0
1
0
0 0 96 782
6 NORMAL
-19 -25 23 -17
4 RLY3
-12 -35 16 -27
2 B1
-5 -45 9 -37
0
17 %D %1 %2 %3 %I %S
0
15 alias:XCONTACTS
4 SIP3
7

0 1 2 3 1 2 3 0
88 0 0 0 1 0 -3 0
3 RLY
4718 0 0
0
0
7 Ground~
168 242 113 0 1 3
0 3
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3874 0 0
0
0
7 Ground~
168 185 113 0 1 3
0 3
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
7 Buffer~
58 148 248 0 2 22
0 20 7
0
0 0 96 90
4 4050
-14 -19 14 -11
3 U2A
13 -5 34 3
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 1 0
1 U
3789 0 0
0
0
11 Contacts:B~
215 155 109 0 10 18
0 11 16 3 0 0 0 0 0 0
1
0
0 0 96 782
6 NORMAL
-19 -25 23 -17
4 RLY1
-12 -35 16 -27
2 B0
-5 -45 9 -37
0
17 %D %1 %2 %3 %I %S
0
15 alias:XCONTACTS
4 SIP3
7

0 1 2 3 1 2 3 0
88 0 0 0 1 0 -2 0
3 RLY
4871 0 0
0
0
7 Op Amp~
219 402 183 0 3 7
0 3 21 2
0
0 0 64 0
5 IDEAL
-18 -25 17 -17
2 U1
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 1 0 0 0
1 U
3750 0 0
0
0
9 Solenoid~
210 148 214 0 10 18
0 7 15 0 0 0 0 0 0 0
1
0
0 0 4192 90
6 5VCOIL
10 0 52 8
4 RLY9
17 -10 45 -2
2 B0
-7 -50 7 -42
0
23 *p=1 r=1
%D %1 0 %I %S
0
11 alias:XCOIL
4 SIP2
5

0 1 2 1 2 0
88 0 0 0 1 0 -2 0
3 RLY
8778 0 0
0
0
9 Solenoid~
210 205 214 0 10 18
0 6 14 0 0 0 0 0 0 0
1
0
0 0 4192 90
6 5VCOIL
10 0 52 8
4 RLY2
17 -10 45 -2
2 B1
-7 -50 7 -42
0
23 *p=1 r=1
%D %1 0 %I %S
0
11 alias:XCOIL
4 SIP2
5

0 1 2 1 2 0
88 0 0 0 1 0 -3 0
3 RLY
538 0 0
0
0
9 Solenoid~
210 262 214 0 10 18
0 5 13 0 0 0 0 0 0 0
1
0
0 0 4192 90
6 5VCOIL
10 0 52 8
4 RLY6
17 -10 45 -2
2 B2
-7 -50 7 -42
0
23 *p=1 r=1
%D %1 0 %I %S
0
11 alias:XCOIL
4 SIP2
5

0 1 2 1 2 0
88 0 0 0 1 0 -4 0
3 RLY
6843 0 0
0
0
9 Solenoid~
210 320 214 0 10 18
0 4 12 0 0 0 0 0 0 0
1
0
0 0 4192 90
6 5VCOIL
10 0 52 8
4 RLY7
17 -10 45 -2
2 B3
-7 -50 7 -42
0
23 *p=1 r=1
%D %1 0 %I %S
0
11 alias:XCOIL
4 SIP2
5

0 1 2 1 2 0
88 0 0 0 1 0 -5 0
3 RLY
3136 0 0
0
0
9 Resistor~
219 399 137 0 2 5
0 21 2
0
0 0 1120 0
2 2k
-7 -14 7 -6
3 R10
-11 -24 10 -16
2 2R
-6 -14 8 -6
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5950 0 0
0
0
9 Resistor~
219 328 146 0 2 5
0 8 21
0
0 0 1120 270
2 2k
8 0 22 8
2 R9
8 -10 22 -2
2 2R
8 -5 22 3
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5670 0 0
0
0
9 Resistor~
219 271 146 0 2 5
0 9 22
0
0 0 1120 270
2 2k
8 0 22 8
2 R7
8 -10 22 -2
2 2R
8 -5 22 3
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6828 0 0
0
0
9 Resistor~
219 300 177 0 2 5
0 22 21
0
0 0 1120 0
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
1 R
-4 -14 3 -6
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6735 0 0
0
0
9 Resistor~
219 214 146 0 2 5
0 10 23
0
0 0 1120 270
2 2k
8 0 22 8
2 R5
8 -10 22 -2
2 2R
8 -5 22 3
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8365 0 0
0
0
9 Resistor~
219 243 177 0 2 5
0 23 22
0
0 0 1120 0
2 1k
-7 -14 7 -6
2 R4
-7 -24 7 -16
1 R
-4 -14 3 -6
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4132 0 0
0
0
9 Resistor~
219 186 177 0 2 5
0 24 23
0
0 0 1120 0
2 1k
-7 -14 7 -6
2 R3
-7 -24 7 -16
1 R
-4 -14 3 -6
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4551 0 0
0
0
9 Resistor~
219 129 177 0 3 5
0 3 24 -1
0
0 0 1120 0
2 2k
-7 -14 7 -6
2 R2
-7 -24 7 -16
2 2R
-7 -14 7 -6
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3635 0 0
0
0
9 Resistor~
219 157 146 0 2 5
0 11 24
0
0 0 1120 270
2 2k
8 0 22 8
2 R1
8 -10 22 -2
2 2R
8 -5 22 3
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3973 0 0
0
0
37
1 2 4 0 0 4224 0 25 5 0 0 2
320 234
320 233
1 2 5 0 0 4224 0 24 6 0 0 2
262 234
262 233
1 2 6 0 0 4224 0 23 7 0 0 2
205 234
205 233
1 2 7 0 0 4224 0 22 19 0 0 2
148 234
148 233
1 1 8 0 0 4224 0 12 27 0 0 2
328 126
328 128
1 1 9 0 0 4224 0 14 28 0 0 2
271 126
271 128
1 1 10 0 0 4224 0 16 30 0 0 2
214 126
214 128
1 1 11 0 0 4224 0 20 34 0 0 2
157 125
157 128
2 0 12 0 0 4480 0 25 0 0 0 3
320 194
320 107
325 107
2 0 13 0 0 4480 0 24 0 0 0 3
262 194
262 107
268 107
2 0 14 0 0 4480 0 23 0 0 0 3
205 194
205 107
211 107
2 0 15 0 0 4480 0 22 0 0 0 3
148 194
148 107
154 107
2 0 16 0 0 4096 0 14 0 0 29 2
256 98
256 83
2 0 16 0 0 0 0 16 0 0 29 2
199 98
199 83
2 0 16 0 0 0 0 20 0 0 29 2
142 97
142 83
3 1 3 0 0 4096 0 20 18 0 0 3
172 97
185 97
185 107
3 1 3 0 0 0 0 16 17 0 0 3
229 98
242 98
242 107
3 1 3 0 0 0 0 14 15 0 0 3
286 98
299 98
299 107
3 1 3 0 0 0 0 12 13 0 0 3
343 98
356 98
356 107
1 1 17 0 0 4224 0 5 1 0 0 2
320 263
320 262
1 1 18 0 0 4224 0 6 2 0 0 2
262 263
262 261
1 1 19 0 0 4224 0 7 3 0 0 2
205 263
205 262
1 1 20 0 0 0 0 19 4 0 0 2
148 263
148 263
1 1 3 0 0 8320 0 9 21 0 0 3
364 202
364 189
384 189
2 0 2 0 0 8320 0 26 0 0 27 3
417 137
436 137
436 183
1 0 21 0 0 8192 0 26 0 0 28 3
381 137
364 137
364 177
3 1 2 0 0 0 0 21 8 0 0 2
420 183
465 183
2 2 21 0 0 4224 0 21 29 0 0 2
384 177
318 177
1 2 16 0 0 4224 0 10 12 0 0 3
113 83
313 83
313 98
1 1 3 0 0 0 0 11 33 0 0 3
103 186
103 177
111 177
2 0 21 0 0 0 0 27 0 0 28 2
328 164
328 177
2 0 22 0 0 4096 0 28 0 0 33 2
271 164
271 177
2 1 22 0 0 4224 0 31 29 0 0 2
261 177
282 177
2 0 23 0 0 4096 0 30 0 0 35 2
214 164
214 177
2 1 23 0 0 4224 0 32 31 0 0 2
204 177
225 177
2 0 24 0 0 4096 0 34 0 0 37 2
157 164
157 177
2 1 24 0 0 4224 0 33 32 0 0 2
147 177
168 177
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
152 324 336 348
156 328 332 344
22 Basic R/2R ladder DAC.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
479 217 521 237
483 221 518 235
5 _____
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
478 216 520 253
482 220 517 248
10 -VREF
  8
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 16
430 223 549 243
434 227 546 241
16 VOUT =       x B
0
1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
572655678 1210432 100 100 0 0
77 66 587 216
7 94 168 164
587 66
77 66
587 66
587 216
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 3e-010 2
1
450 183
0 2 0 0 1	0 27 0 0
829752294 8550464 100 100 0 0
77 66 587 246
4 405 625 740
586 66
77 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 1e-006 10
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
