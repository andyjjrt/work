CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 460
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 460
10485778 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 133 233 0 1 11
0 18
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
13 D (Direction)
-106 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
2 +V
167 593 86 0 1 3
0 3
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
14 Logic Display~
6 298 27 0 1 2
10 9
0
0 0 54384 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
1 B
-4 -21 3 -13
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 317 27 0 1 2
10 10
0
0 0 54384 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
1 A
-4 -21 3 -13
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
2 +V
167 270 95 0 1 3
0 13
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
2 +V
167 109 95 0 1 3
0 14
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
9 Inverter~
13 216 116 0 2 22
0 19 20
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
9914 0 0
0
0
7 Pulser~
4 46 195 0 10 12
0 21 22 17 23 0 0 5 5 6
7
0
0 0 5168 0
0
2 V2
-7 -28 7 -20
4 Step
-14 -28 14 -20
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3747 0 0
0
0
9 2-In XOR~
219 330 138 0 3 22
0 10 18 15
0
0 0 112 0
6 74LS86
-21 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 2 3 0
1 U
3549 0 0
0
0
9 2-In XOR~
219 176 157 0 3 22
0 9 18 19
0
0 0 112 0
6 74LS86
-21 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0
65 0 0 0 4 1 3 0
1 U
7931 0 0
0
0
9 Inverter~
13 44 148 0 2 22
0 15 16
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
9325 0 0
0
0
6 74113~
219 270 146 0 6 22
0 20 17 19 13 12 10
0
0 0 4208 0
7 74LS113
-25 -42 24 -34
3 U1B
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 2 1 0
1 U
8903 0 0
0
0
6 74113~
219 109 147 0 6 22
0 15 17 16 14 11 9
0
0 0 4208 0
7 74LS113
-25 -42 24 -34
3 U1A
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 1 1 0
1 U
3834 0 0
0
0
14 Opto Isolator~
173 448 89 0 64 64
0 10 2 6 2 0 0 0 0 0
10 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162722
0
0 0 112 0
7 OPTOISO
-26 -28 23 -20
2 U7
-9 -38 5 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
5

0 1 2 3 4 0
88 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
14 Opto Isolator~
173 448 125 0 64 64
0 12 2 7 2 0 0 0 0 0
10 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162720
0
0 0 112 0
7 OPTOISO
-26 -28 23 -20
2 U6
-9 -38 5 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
5

0 1 2 3 4 0
88 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
14 Opto Isolator~
173 448 161 0 64 64
0 9 2 5 2 0 0 0 0 0
10 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162720
0
0 0 112 0
7 OPTOISO
-26 -28 23 -20
2 U5
-9 -38 5 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
5

0 1 2 3 4 0
88 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
14 Opto Isolator~
173 448 197 0 64 64
0 11 2 4 2 0 0 0 0 0
10 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 2162694
0
0 0 112 0
7 OPTOISO
-26 -28 23 -20
2 U4
-9 -38 5 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
5

0 1 2 3 4 0
88 0 0 0 1 0 0 0
1 U
3874 0 0
0
0
7 Ground~
168 481 232 0 1 3
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6671 0 0
0
0
8 Stepper~
185 550 131 0 6 13
13 6 3 7 5 3 4
0
0 0 4208 0
4 100H
10 -16 38 -8
2 M1
17 -26 31 -18
0
0
130 %DA %1 N%DA %V
R%DA N%DA %2 10
%DB %3 N%DB %V
R%DB N%DB %2 10
%DC %4 N%DC %V
R%DC N%DC %5 10
%DD %6 N%DD %V
R%DD N%DD %5 10
0
0
4 SIP6
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
76 0 0 0 1 1 0 0
1 M
3789 0 0
0
0
35
2 0 3 0 0 4096 0 19 0 0 13 2
586 107
593 107
3 6 4 0 0 4224 0 17 19 0 0 4
474 185
511 185
511 161
514 161
3 4 5 0 0 4224 0 16 19 0 0 2
474 149
514 149
3 1 6 0 0 4224 0 14 19 0 0 4
474 77
511 77
511 101
514 101
3 3 7 0 0 4224 0 15 19 0 0 2
474 113
514 113
0 0 8 0 0 4480 0 0 0 0 0 5
397 52
397 251
501 251
501 52
399 52
1 0 9 0 0 4096 0 3 0 0 10 2
298 45
298 61
1 0 10 0 0 4096 0 4 0 0 12 2
317 45
317 77
5 1 11 0 0 12416 0 13 17 0 0 6
139 148
146 148
146 69
375 69
375 185
420 185
0 1 9 0 0 8320 0 0 16 31 0 5
152 130
152 61
382 61
382 149
420 149
5 1 12 0 0 8320 0 12 15 0 0 3
300 147
300 113
420 113
0 1 10 0 0 8320 0 0 14 35 0 3
308 129
308 77
420 77
1 5 3 0 0 4224 0 2 19 0 0 3
593 95
593 155
586 155
2 0 2 0 0 4096 0 17 0 0 17 2
420 209
412 209
2 0 2 0 0 0 0 16 0 0 17 2
420 173
412 173
2 0 2 0 0 0 0 15 0 0 17 2
420 137
412 137
2 0 2 0 0 8320 0 14 0 0 21 4
420 101
412 101
412 226
481 226
4 0 2 0 0 0 0 15 0 0 21 2
474 137
481 137
4 0 2 0 0 0 0 16 0 0 21 2
474 173
481 173
4 0 2 0 0 0 0 17 0 0 21 2
474 209
481 209
4 1 2 0 0 0 0 14 18 0 0 3
474 101
481 101
481 226
1 4 13 0 0 4224 0 5 12 0 0 2
270 104
270 102
1 4 14 0 0 4224 0 6 13 0 0 2
109 104
109 103
1 0 15 0 0 8192 0 13 0 0 25 3
85 130
78 130
78 53
3 1 15 0 0 12416 0 9 11 0 0 5
363 138
367 138
367 53
29 53
29 148
2 3 16 0 0 4224 0 11 13 0 0 2
65 148
85 148
2 0 17 0 0 4096 0 13 0 0 28 2
78 139
78 186
3 2 17 0 0 4224 0 8 12 0 0 3
70 186
239 186
239 138
2 0 18 0 0 8192 0 10 0 0 30 3
160 166
152 166
152 233
1 2 18 0 0 4224 0 1 9 0 0 4
145 233
308 233
308 147
314 147
6 1 9 0 0 0 0 13 10 0 0 4
133 130
152 130
152 148
160 148
0 1 19 0 0 4224 0 0 7 33 0 5
220 157
220 130
193 130
193 116
201 116
3 3 19 0 0 0 0 10 12 0 0 4
209 157
231 157
231 147
246 147
2 1 20 0 0 4224 0 7 12 0 0 3
237 116
237 129
246 129
6 1 10 0 0 0 0 12 9 0 0 2
294 129
314 129
2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 206
25 283 585 347
29 287 581 335
206 A synchronous counter supplies the appropriate sequential outputs 
to drive a stepper motor. (Note: In this configuration, the stepper 
runs in the opposite direction from the one described in the text.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 21
394 18 478 55
398 22 475 50
21 Current 
amplifiers
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
