CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 8 100 9
4 70 635 440
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 440 635 571
27262994 0
0
6 Title:
5 Name:
0
0
0
14
14 Logic Display~
6 470 30 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8953 0 0
0
0
14 Logic Display~
6 354 31 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 234 31 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
6 74113~
219 188 130 0 6 22
0 8 3 8 8 10 4
0
0 0 4192 0
7 74LS113
-25 -42 24 -34
3 U1A
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 1 0
1 U
6153 0 0
0
0
6 74113~
219 298 130 0 6 22
0 7 2 7 7 11 3
0
0 0 4192 0
7 74LS113
-25 -42 24 -34
3 U1B
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 2 1 0
1 U
5394 0 0
0
0
6 74113~
219 411 130 0 6 22
0 6 5 6 6 12 2
0
0 0 4192 0
7 74LS113
-25 -42 24 -34
3 U2A
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 2 0
1 U
7734 0 0
0
0
2 +V
167 150 75 0 1 3
0 8
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
2 +V
167 259 75 0 1 3
0 7
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
2 +V
167 371 78 0 1 3
0 6
0
0 0 53472 0
2 5V
-7 -22 7 -14
3 V10
-11 -32 10 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3549 0 0
0
0
7 Pulser~
4 272 212 0 10 12
0 13 14 5 15 0 0 10 10 11
7
0
0 0 4128 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7931 0 0
0
0
5 SCOPE
12 331 192 0 1 11
0 5
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
5 SCOPE
12 447 36 0 1 11
0 2
0
0 0 57568 0
2 Q0
-8 -4 6 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
5 SCOPE
12 331 37 0 1 11
0 3
0
0 0 57568 0
2 Q1
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
5 SCOPE
12 211 37 0 1 11
0 4
0
0 0 57568 0
2 Q2
-8 -4 6 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
21
0 0 9 0 0 16 0 0 0 0 0 5
310 266
581 266
581 299
310 299
310 266
1 0 2 0 0 4096 0 1 0 0 6 2
470 48
447 48
1 0 3 0 0 4096 0 2 0 0 7 2
354 49
331 49
1 0 4 0 0 4096 0 3 0 0 8 2
234 49
211 49
1 0 5 0 0 4096 0 11 0 0 19 2
331 204
331 203
1 0 2 0 0 4096 0 12 0 0 18 2
447 48
447 113
1 0 3 0 0 0 0 13 0 0 20 2
331 49
331 56
1 6 4 0 0 4224 0 14 4 0 0 3
211 49
211 113
212 113
1 0 6 0 0 4096 0 6 0 0 10 2
387 113
371 113
3 0 6 0 0 8320 0 6 0 0 15 3
387 131
371 131
371 87
1 0 7 0 0 4096 0 5 0 0 12 2
274 113
259 113
0 3 7 0 0 4224 0 0 5 16 0 3
259 86
259 131
274 131
1 0 8 0 0 4096 0 4 0 0 14 2
164 113
150 113
0 3 8 0 0 4224 0 0 4 17 0 3
150 86
150 131
164 131
1 4 6 0 0 0 0 9 6 0 0 3
371 87
411 87
411 86
1 4 7 0 0 0 0 8 5 0 0 3
259 84
259 86
298 86
1 4 8 0 0 0 0 7 4 0 0 3
150 84
150 86
188 86
6 2 2 0 0 12416 0 6 5 0 0 6
435 113
447 113
447 169
249 169
249 122
267 122
2 3 5 0 0 8320 0 6 10 0 0 4
380 122
362 122
362 203
296 203
6 2 3 0 0 12416 0 5 4 0 0 6
322 113
331 113
331 56
126 56
126 122
157 122
0 6 2 0 0 0 0 0 6 18 0 2
435 113
435 113
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
312 263 578 300
316 267 575 295
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 3
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 65
27 256 219 320
31 260 215 308
65 J-K flip-flops wired 
as a three-bit binary 
counter (MOD-8).
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
