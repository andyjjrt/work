CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 21 100 9
4 70 635 393
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 393
8388626 0
0
6 Title:
5 Name:
0
0
0
6
13 Logic Switch~
5 83 131 0 1 11
0 4
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
5 CLEAR
-54 -5 -19 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 83 47 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21616 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
3 SET
-39 -4 -18 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
14 Logic Display~
6 230 97 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 230 32 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
5 4011~
219 152 122 0 3 22
0 2 4 3
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
5394 0 0
0
0
5 4011~
219 152 56 0 3 22
0 5 3 2
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
7734 0 0
0
0
10
0 1 2 0 0 8336 0 0 5 4 0 5
184 56
184 82
124 82
124 113
128 113
2 0 3 0 0 12416 0 6 0 0 3 5
128 65
110 65
110 96
185 96
185 122
1 3 3 0 0 0 0 3 5 0 0 3
230 115
230 122
179 122
1 3 2 0 0 0 0 4 6 0 0 3
230 50
230 56
179 56
2 1 4 0 0 4224 0 5 1 0 0 2
128 131
95 131
1 1 5 0 0 4224 0 6 2 0 0 2
128 47
95 47
0 0 1 0 0 4256 0 0 0 0 0 2
428 35
428 117
0 0 6 0 0 4224 0 0 0 0 0 2
338 117
510 117
0 0 7 0 0 4224 0 0 0 0 0 2
338 50
510 50
0 0 8 0 0 4224 0 0 0 0 0 2
338 35
510 35
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
233 108 249 132
237 112 245 128
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
233 100 249 124
237 104 245 120
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
135 163 167 187
139 167 163 183
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
407 163 439 187
411 167 435 183
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 117
337 31 521 175
341 35 517 147
117 Set  Clear   Output
 1     1    No change
 0     1    Q=1
 1     0    Q=0
 0     0    Invalid*

*produces Q=Q=1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
433 119 449 143
437 123 445 139
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 31
210 207 346 251
214 211 342 243
31 (a) NAND latch
(b) truth table
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
231 43 247 67
235 47 243 63
1 Q
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 2e-005 1e-008 1e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
