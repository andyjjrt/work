CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 430
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 430 635 754
25165842 0
0
6 Title:
5 Name:
0
0
0
16
5 74147
219 392 149 0 13 27
0 6 7 8 9 10 11 12 13 14
2 3 4 5
0
0 0 12512 0
5 74147
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
121 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
27

0 10 5 4 3 2 1 13 12 11
9 7 6 14 10 5 4 3 2 1
13 12 11 9 7 6 14 0
65 0 0 0 1 0 0 0
1 U
8953 0 0
0
0
9 Data Seq~
170 114 149 0 17 18
0 7 8 9 10 11 12 13 14 16
17 1 1 20 20 21 0 33
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
4441 0 0
0
0
AAPPAAAAIAMAOAPAPIPMPOAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
9 Data Seq~
170 114 71 0 17 18
0 18 19 20 21 22 23 24 6 25
26 1 1 20 20 21 0 33
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS2
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
3618 0 0
0
0
AAABAAABABABABABABABABAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA
5 SCOPE
12 174 79 0 1 11
0 14
0
0 0 57568 0
3 A1n
-11 -4 10 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
5 SCOPE
12 195 93 0 1 11
0 13
0
0 0 57568 0
3 A2n
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 215 79 0 1 11
0 12
0
0 0 57568 0
3 A3n
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 235 93 0 1 11
0 11
0
0 0 57568 0
3 A4n
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 255 79 0 1 11
0 10
0
0 0 57568 0
3 A5n
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 275 93 0 1 11
0 9
0
0 0 57568 0
3 A6n
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 295 79 0 1 11
0 8
0
0 0 57568 0
3 A7n
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
5 SCOPE
12 315 93 0 1 11
0 7
0
0 0 57568 0
3 A8n
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
5 SCOPE
12 335 79 0 1 11
0 6
0
0 0 57568 0
3 A9n
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
5 SCOPE
12 507 113 0 1 11
0 2
0
0 0 57568 0
3 O0n
-11 -4 10 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
5 SCOPE
12 487 99 0 1 11
0 3
0
0 0 57568 0
3 O1n
-10 -4 11 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
5 SCOPE
12 467 113 0 1 11
0 4
0
0 0 57568 0
3 O2n
-10 -4 11 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7668 0 0
0
0
5 SCOPE
12 446 99 0 1 11
0 5
0
0 0 57568 0
3 O3n
-10 -4 11 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4718 0 0
0
0
23
0 0 15 0 0 16 0 0 0 0 0 5
315 246
586 246
586 279
315 279
315 246
10 1 2 0 0 4224 0 1 13 0 0 3
430 158
507 158
507 125
11 1 3 0 0 4224 0 1 14 0 0 3
430 149
487 149
487 111
12 1 4 0 0 4224 0 1 15 0 0 3
430 140
467 140
467 125
13 1 5 0 0 8320 0 1 16 0 0 3
430 131
446 131
446 111
1 0 6 0 0 4096 0 12 0 0 15 2
335 91
335 113
1 0 7 0 0 4096 0 11 0 0 16 2
315 105
315 122
1 0 8 0 0 4096 0 10 0 0 17 2
295 91
295 131
1 0 9 0 0 4096 0 9 0 0 18 2
275 105
275 140
1 0 10 0 0 4096 0 8 0 0 19 2
255 91
255 149
1 0 11 0 0 4096 0 7 0 0 20 2
235 105
235 158
1 0 12 0 0 4096 0 6 0 0 21 2
215 91
215 167
1 0 13 0 0 4096 0 5 0 0 22 2
195 105
195 176
1 0 14 0 0 4096 0 4 0 0 23 2
174 91
174 185
8 1 6 0 0 8320 0 3 1 0 0 3
146 107
146 113
354 113
1 2 7 0 0 4224 0 2 1 0 0 2
146 122
354 122
2 3 8 0 0 4224 0 2 1 0 0 2
146 131
354 131
3 4 9 0 0 4224 0 2 1 0 0 2
146 140
354 140
4 5 10 0 0 4224 0 2 1 0 0 2
146 149
354 149
5 6 11 0 0 4224 0 2 1 0 0 2
146 158
354 158
6 7 12 0 0 4224 0 2 1 0 0 2
146 167
354 167
7 8 13 0 0 4224 0 2 1 0 0 2
146 176
354 176
8 9 14 0 0 4224 0 2 1 0 0 2
146 185
354 185
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
317 243 583 280
321 247 580 275
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 41
44 245 220 289
48 249 216 281
41 74147 decimal-to-BCD 
priority encoder.
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
267780172 8525888 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
9.98039 0 5.4 0 10 10
12401 0
4 1e-006 2
2
221 112
0 7 0 0 2	0 24 0 0
367 106
0 2 0 0 1	0 24 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 24 0 0
200 112
0 7 0 0 2	0 24 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
