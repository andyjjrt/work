CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 432
8388626 0
0
6 Title:
5 Name:
0
0
0
4
13 Logic Switch~
5 302 181 0 1 11
0 3
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
18 Excessive Pressure
-151 -3 -25 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 301 123 0 1 11
0 4
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
21 Excessive Temperature
-172 -5 -25 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
8 2-In OR~
219 365 151 0 3 22
0 4 3 2
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3618 0 0
0
0
14 Logic Display~
6 426 133 0 1 2
10 2
0
0 0 54384 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
5 Alarm
-19 -28 16 -20
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
3
3 1 2 0 0 4224 0 3 4 0 0 2
398 151
426 151
1 2 3 0 0 4224 0 1 3 0 0 4
314 181
344 181
344 160
352 160
1 1 4 0 0 4224 0 2 3 0 0 4
313 123
344 123
344 142
352 142
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 52
76 263 500 287
80 267 496 283
52 Example of the use of an OR gate in an alarm system.
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
