CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 432 635 558
25165842 0
0
6 Title:
5 Name:
0
0
0
7
2 +V
167 233 98 0 1 3
0 3
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8953 0 0
0
0
5 SCOPE
12 118 114 0 1 11
0 7
0
0 0 57568 0
1 J
-4 -4 3 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 153 114 0 1 11
0 6
0
0 0 57568 0
1 K
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 188 114 0 1 11
0 5
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
5 SCOPE
12 275 113 0 1 11
0 4
0
0 0 57568 0
1 Q
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
9 Data Seq~
170 62 116 0 17 18
0 11 12 13 14 15 7 5 6 16
17 33 5 50 5 5 0 51
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
7734 0 0
0
0
AAAAAAACACAAABADAHAFAFAHACAAAAACAGAEAEAGAHAFAFAHAHAFAFAHIHAAAAAAAAAAAAAAAAAAAAAA
AAAAAAAAAAAAAAAAAAAAAA
6 74113~
219 233 151 0 6 22
0 7 5 6 3 18 4
0
0 0 4192 0
6 74F113
-22 -42 20 -34
3 U2A
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 1 5 0
1 U
9914 0 0
0
0
13
1 4 3 0 0 16 0 1 7 0 0 2
233 107
233 107
1 6 4 0 0 16 0 5 7 0 0 3
275 125
275 134
257 134
1 0 5 0 0 16 0 4 0 0 7 2
188 126
188 143
1 0 6 0 0 16 0 3 0 0 6 2
153 126
153 152
1 0 7 0 0 16 0 2 0 0 8 2
118 126
118 134
8 3 6 0 0 16 0 6 7 0 0 2
94 152
209 152
7 2 5 0 0 16 0 6 7 0 0 2
94 143
202 143
6 1 7 0 0 16 0 6 7 0 0 2
94 134
209 134
0 0 1 0 0 48 0 0 0 10 12 2
437 89
437 173
0 0 8 0 0 16 0 0 0 0 0 2
343 89
564 89
0 0 9 0 0 16 0 0 0 0 0 2
343 105
564 105
0 0 10 0 0 16 0 0 0 0 0 2
343 173
564 173
0 0 2 0 0 0 0 0 0 0 0 5
318 261
589 261
589 294
318 294
318 261
15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
405 99 421 123
409 103 417 119
1 |
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
405 103 421 127
409 107 417 123
1 v
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
405 118 421 142
409 122 417 138
1 v
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
405 114 421 138
409 118 417 134
1 |
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
406 133 422 157
410 137 418 153
1 v
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
406 129 422 153
410 133 418 149
1 |
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
406 150 422 174
410 154 418 170
1 v
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
406 146 422 170
410 150 418 166
1 |
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 43
442 86 570 190
446 90 566 170
43       Q
Qo (no change)
1
0
Qo (toggles)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
397 86 429 110
401 90 425 106
3 CLK
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
350 86 374 190
354 90 370 170
13 J
0
1
0
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
377 86 401 190
381 90 397 170
13 K
0
0
1
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
442 136 466 160
446 140 462 156
2 __
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
320 258 586 295
324 262 583 290
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 74
12 256 308 300
16 260 304 292
74 Clocked J-K flip-flop that triggers 
only on negative-going transitions.
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 4.6e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.006 0 5.4 0 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
