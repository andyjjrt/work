CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 436
11010066 0
0
6 Title:
5 Name:
0
0
0
8
9 2-In AND~
219 274 87 0 3 22
0 3 4 7
0
0 0 112 512
6 74LS08
-21 -24 21 -16
3 U2A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8953 0 0
0
0
9 Terminal~
194 405 169 0 1 3
0 2
0
0 0 49520 270
2 Q0
2 -5 16 3
2 T4
-7 -25 7 -17
0
3 Q0;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4441 0 0
0
0
9 Terminal~
194 405 160 0 1 3
0 3
0
0 0 49520 270
2 Q1
2 -5 16 3
2 T3
-7 -25 7 -17
0
3 Q1;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3618 0 0
0
0
9 Terminal~
194 405 151 0 1 3
0 4
0
0 0 49520 270
2 Q2
2 -5 16 3
2 T2
-7 -25 7 -17
0
3 Q2;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
6153 0 0
0
0
9 Terminal~
194 440 142 0 1 3
0 5
0
0 0 49520 270
2 Q3
2 -5 16 3
2 T1
-7 -25 7 -17
0
3 Q3;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
5394 0 0
0
0
7 Ground~
168 169 177 0 1 3
0 6
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
11 Signal Gen~
195 128 164 0 24 64
0 8 6 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1176256512 0 1084227584
944879383 897988541 897988541 944879383 953267991
20
0 10000 0 5 5e-005 1e-006 1e-006 5e-005 0.0001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 80 0
4 0/5V
-15 -30 13 -22
2 V2
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 PULSE(0 5 50u 1u 1u 50u 100u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
7 74LS293
154 275 150 0 8 17
0 7 5 8 2 5 4 3 2
0
0 0 12528 0
7 74LS293
-24 -35 25 -27
2 U1
-7 -36 7 -28
0
15 DVCC=14;DGND=7;
77 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP14
17

0 12 13 10 11 8 4 5 9 12
13 10 11 8 4 5 9 0
65 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
11
3 1 7 0 0 8320 0 1 8 0 0 4
249 87
221 87
221 141
243 141
1 0 3 0 0 8208 0 1 0 0 5 3
294 78
339 78
339 159
2 0 4 0 0 8192 0 1 0 0 6 3
294 96
328 96
328 150
0 2 5 0 0 8192 0 0 8 7 0 5
317 141
317 113
231 113
231 150
243 150
1 7 3 0 0 4224 0 3 8 0 0 2
393 159
307 159
1 6 4 0 0 4224 0 4 8 0 0 2
393 150
307 150
1 5 5 0 0 4224 0 5 8 0 0 2
428 141
307 141
1 8 2 0 0 4096 0 2 8 0 0 2
393 168
307 168
1 2 6 0 0 8320 0 6 7 0 0 3
169 171
169 169
159 169
1 3 8 0 0 4224 0 7 8 0 0 2
159 159
237 159
0 4 2 0 0 8320 0 0 8 8 0 5
318 168
318 187
231 187
231 168
237 168
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 20
436 115 583 135
440 119 580 133
20 f = 10kHz/14 = 714Hz
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 74
139 269 451 313
143 273 447 305
74 An external AND gate is needed to 
wire the 74LS293 as a MOD-14 counter.
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.003 6e-006 6e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
62522106 8550464 100 100 0 0
77 66 587 246
3 436 635 771
451 66
213 66
587 66
587 246
0 0
0.0022 0.0008 30 -30 0.003 0.003
13425 0
2 0.0005 10
5
182 159
0 8 0 60 1	0 10 0 0
385 141
0 5 0 -59 1	0 7 0 0
375 150
0 4 0 -29 1	0 6 0 0
363 159
0 3 0 0 1	0 5 0 0
352 168
0 2 0 32 1	0 8 0 0
110889084 8550464 100 100 0 0
77 66 587 246
3 436 635 771
442 66
170 66
587 66
587 182
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 0.001 2
1
348 141
0 4 0 0 1	0 5 0 0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
