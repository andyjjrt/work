CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 1 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 432
8388626 0
0
6 Title:
5 Name:
0
0
0
9
7 74LS191
135 175 173 0 14 29
0 2 7 8 2 2 2 2 2 10
11 6 5 4 3
0
0 0 12512 0
7 74LS191
-24 -51 25 -43
2 U1
-7 -52 7 -44
0
15 DVCC=16;DGND=8;
122 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 4 14 11 5 9 10 1 15 13
12 7 6 2 3 4 14 11 5 9
10 1 15 13 12 7 6 2 3 0
65 0 0 512 1 0 0 0
1 U
8953 0 0
0
0
2 +V
167 117 126 0 1 3
0 8
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 126 236 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Pulser~
4 61 164 0 10 12
0 12 13 7 14 0 0 5 5 6
7
0
0 0 4128 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
6153 0 0
0
0
12 Hex Display~
7 302 148 0 16 19
10 3 4 5 6 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5394 0 0
0
0
14 Logic Display~
6 225 140 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 236 140 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 247 140 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 258 140 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
17
1 0 3 0 0 4096 0 9 0 0 5 2
258 158
258 209
1 0 4 0 0 4096 0 8 0 0 6 2
247 158
247 200
1 0 5 0 0 4096 0 7 0 0 7 2
236 158
236 191
1 0 6 0 0 4096 0 6 0 0 8 2
225 158
225 182
1 14 3 0 0 8320 0 5 1 0 0 3
311 172
311 209
207 209
2 13 4 0 0 8320 0 5 1 0 0 3
305 172
305 200
207 200
3 12 5 0 0 8320 0 5 1 0 0 3
299 172
299 191
207 191
4 11 6 0 0 8320 0 5 1 0 0 3
293 172
293 182
207 182
8 0 2 0 0 4096 0 1 0 0 15 2
143 209
126 209
7 0 2 0 0 0 0 1 0 0 15 2
143 200
126 200
6 0 2 0 0 0 0 1 0 0 15 2
143 191
126 191
5 0 2 0 0 0 0 1 0 0 15 2
143 182
126 182
4 0 2 0 0 0 0 1 0 0 15 2
143 173
126 173
3 2 7 0 0 4224 0 4 1 0 0 2
85 155
143 155
1 1 2 0 0 8320 0 1 3 0 0 3
137 146
126 146
126 230
1 3 8 0 0 4224 0 2 1 0 0 3
117 135
117 164
137 164
0 0 9 0 0 4224 0 0 0 0 0 2
339 34
584 34
6
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 41
9 272 225 316
13 276 221 308
41 Hexadecimal number system 
and counter.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
213 97 269 121
217 101 265 117
6 Binary
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
287 97 319 121
291 101 315 117
3 Hex
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 123
341 15 437 359
345 19 433 291
123 Hexadecimal
    0
    1
    2
    3
    4
    5
    6
    7
    8
    9
    A
    B
    C
    D
    E
    F
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 103
451 16 515 360
455 20 511 292
103 Decimal
   0
   1
   2
   3
   4
   5
   6
   7
   8
   9
  10
  11
  12
  13
  14
  15
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 118
527 15 583 359
531 19 579 291
118 Binary
 0000
 0001
 0010
 0011
 0100
 0101
 0110
 0111
 1000
 1001
 1010
 1011
 1100
 1101
 1110
 1111
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
