CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 563
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 563
8912918 0
0
6 Title:
5 Name:
0
0
0
19
13 Logic Switch~
5 182 290 0 1 11
0 8
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 B
-29 -3 -22 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 181 209 0 1 11
0 7
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 A
-28 -3 -21 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
9 Terminal~
194 400 227 0 1 3
0 2
0
0 0 49520 270
1 X
-7 -14 0 -6
2 T1
3 -17 17 -9
0
2 X;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
3618 0 0
0
0
7 Ground~
168 433 238 0 1 3
0 3
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
11 Multimeter~
205 408 187 0 21 21
0 2 15 16 3 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
7 Ground~
168 344 328 0 1 3
0 3
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
2 +V
167 321 95 0 1 3
0 9
0
0 0 53616 0
3 +5V
-10 -15 11 -7
2 V1
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
12 NPN Trans:B~
219 339 252 0 3 7
0 2 4 3
0
0 0 592 0
6 2N2270
7 0 49 8
2 Q6
2 -3 16 5
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3747 0 0
0
0
6 Diode~
219 344 208 0 2 5
0 13 2
0
0 0 592 270
5 DIODE
11 0 46 8
2 D1
12 -5 26 3
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3549 0 0
0
0
12 NPN Trans:B~
219 339 176 0 3 7
0 14 5 13
0
0 0 592 0
6 2N2270
7 0 49 8
2 Q5
2 -3 16 5
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
7931 0 0
0
0
12 NPN Trans:B~
219 275 209 0 3 7
0 5 10 4
0
0 0 592 0
6 2N2270
7 0 49 8
2 Q3
3 -3 17 5
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
9325 0 0
0
0
12 NPN Trans:B~
219 231 202 0 3 7
0 10 12 7
0
0 0 592 270
6 2N2270
-23 30 19 38
2 Q1
-7 6 7 14
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
8903 0 0
0
0
12 NPN Trans:B~
219 232 283 0 3 7
0 6 11 8
0
0 0 592 270
6 2N2270
-23 30 19 38
2 Q2
-8 7 6 15
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3834 0 0
0
0
12 NPN Trans:B~
219 269 290 0 3 7
0 5 6 4
0
0 0 592 0
6 2N2270
7 0 49 8
2 Q4
2 -4 16 4
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-39
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3363 0 0
0
0
9 Resistor~
219 344 134 0 3 5
0 9 14 1
0
0 0 880 270
3 130
7 0 28 8
2 R4
10 -10 24 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7668 0 0
0
0
9 Resistor~
219 298 134 0 3 5
0 9 5 1
0
0 0 880 270
4 1.6k
8 0 36 8
2 R3
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4718 0 0
0
0
9 Resistor~
219 229 137 0 3 5
0 9 12 1
0
0 0 880 270
2 4k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
9 Resistor~
219 230 247 0 3 5
0 9 11 1
0
0 0 880 270
2 4k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6671 0 0
0
0
9 Resistor~
219 319 313 0 4 5
0 4 3 0 -1
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3789 0 0
0
0
24
0 3 4 0 0 4240 0 0 11 5 0 3
288 313
288 227
280 227
1 0 5 0 0 12432 0 14 0 0 20 4
274 272
274 269
298 269
298 176
1 2 6 0 0 4240 0 13 14 0 0 2
248 290
251 290
2 0 3 0 0 4112 0 19 0 0 6 2
337 313
344 313
3 1 4 0 0 16 0 14 19 0 0 3
274 308
274 313
301 313
1 3 3 0 0 4240 0 6 8 0 0 2
344 322
344 270
3 1 7 0 0 4240 0 12 2 0 0 2
211 209
193 209
3 1 8 0 0 4240 0 13 1 0 0 2
212 290
194 290
1 0 9 0 0 12432 0 18 0 0 18 4
230 229
230 225
255 225
255 109
1 2 10 0 0 4240 0 12 11 0 0 4
247 209
258 209
258 209
257 209
2 2 11 0 0 4240 0 18 13 0 0 2
230 265
230 267
2 2 12 0 0 4240 0 17 12 0 0 2
229 155
229 186
1 0 2 0 0 4112 0 5 0 0 14 2
383 210
383 226
0 1 2 0 0 4240 0 0 3 21 0 2
344 226
388 226
1 0 9 0 0 16 0 7 0 0 18 2
321 104
321 109
1 4 3 0 0 16 0 4 5 0 0 2
433 232
433 210
1 0 9 0 0 16 0 16 0 0 18 2
298 116
298 109
1 1 9 0 0 16 0 17 15 0 0 4
229 119
229 109
344 109
344 116
2 0 4 0 0 16 0 8 0 0 1 2
321 252
288 252
2 0 5 0 0 16 0 10 0 0 24 3
321 176
298 176
298 162
2 1 2 0 0 16 0 9 8 0 0 2
344 218
344 234
3 1 13 0 0 4240 0 10 9 0 0 2
344 194
344 198
2 1 14 0 0 4240 0 15 10 0 0 2
344 152
344 158
2 1 5 0 0 16 0 16 11 0 0 4
298 152
298 162
280 162
280 191
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
205 404 381 428
209 408 377 424
21 TTL NOR gate circuit.
22 .OPTIONS RSHUNT=1E12

1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
160958526 1210432 100 100 0 0
77 66 587 216
8 92 169 162
587 66
77 66
587 66
587 216
0 0
0.016 0 24 0 0.016 24
12401 0
4 2 2
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
