CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 432
8388626 0
0
6 Title:
5 Name:
0
0
0
4
13 Logic Switch~
5 331 133 0 1 11
0 3
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 B
-22 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 331 95 0 1 11
0 4
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-22 -1 -15 7
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 458 95 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
8 2-In OR~
219 386 114 0 3 22
0 4 3 2
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6153 0 0
0
0
7
0 0 1 0 0 4256 0 0 0 0 0 2
165 76
165 158
1 3 2 0 0 8320 0 3 4 0 0 3
458 113
458 114
419 114
2 1 3 0 0 12416 0 4 1 0 0 4
373 123
359 123
359 133
343 133
1 1 4 0 0 12416 0 4 2 0 0 4
373 105
359 105
359 95
343 95
0 0 5 0 0 4224 0 0 0 0 0 2
107 158
219 158
0 0 6 0 0 4224 0 0 0 0 0 2
107 76
218 76
0 0 7 0 0 4224 0 0 0 0 0 2
107 92
219 92
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 74
109 248 453 292
113 252 449 284
74 (a) Truth table defining the OR operation;
(b) two-input OR gate circuit.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
171 72 219 176
175 76 215 156
25 x=A+B
  0
  1
  1
  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
138 72 162 176
142 76 158 156
13 B
0
1
0
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
111 72 135 176
115 76 131 156
13 A
0
0
1
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
152 54 176 78
156 58 172 74
2 OR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
147 179 179 203
151 183 175 199
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
433 117 481 141
437 121 477 137
5 x=A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
366 187 398 211
370 191 394 207
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
354 171 418 195
358 175 414 191
7 OR Gate
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
