CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 426
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 426
8388626 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 71 63 0 1 11
0 10
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 D
-23 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 72 114 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 22128 0
2 5V
-6 -16 8 -8
6 ENABLE
-57 -9 -15 -1
4 (EN)
-49 1 -21 9
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
5 4011~
219 175 72 0 3 22
0 10 11 8
0
0 0 1136 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
1 1
-8 -4 -1 4
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
3618 0 0
0
0
5 4011~
219 175 158 0 3 22
0 11 9 7
0
0 0 1136 0
4 4011
-7 -24 21 -16
3 U1B
-12 -25 9 -17
1 2
-7 -4 0 4
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 1 0
1 U
6153 0 0
0
0
13 2-In NAND:DM~
219 267 81 0 3 22
0 8 6 5
0
0 0 1136 0
4 4011
-7 -24 21 -16
3 U2A
-3 -25 18 -17
1 3
4 -4 11 4
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 2 0
1 U
5394 0 0
0
0
13 2-In NAND:DM~
219 268 149 0 3 22
0 5 7 6
0
0 0 1136 0
4 4011
-7 -24 21 -16
3 U2B
-3 -25 18 -17
1 4
4 -4 11 4
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
7734 0 0
0
0
9 Inverter~
13 121 167 0 2 22
0 10 9
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
9914 0 0
0
0
14 Logic Display~
6 337 60 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 337 128 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
15
0 0 1 0 0 4272 0 0 0 0 0 2
447 49
447 115
0 0 2 0 0 4240 0 0 0 0 0 2
383 115
571 115
0 0 3 0 0 4240 0 0 0 0 0 2
383 64
571 64
0 0 4 0 0 4240 0 0 0 0 0 2
383 49
571 49
0 1 5 0 0 8320 0 0 6 8 0 5
307 81
307 107
250 107
250 140
249 140
2 0 6 0 0 12416 0 5 0 0 7 5
248 90
240 90
240 122
307 122
307 149
1 3 6 0 0 0 0 9 6 0 0 5
337 146
337 149
298 149
298 149
301 149
1 3 5 0 0 0 0 8 5 0 0 3
337 78
337 81
300 81
2 3 7 0 0 4224 0 6 4 0 0 2
249 158
202 158
1 3 8 0 0 4224 0 5 3 0 0 2
248 72
202 72
2 2 9 0 0 4224 0 4 7 0 0 2
151 167
142 167
0 1 10 0 0 4224 0 0 7 13 0 3
97 63
97 167
106 167
1 1 10 0 0 0 0 3 1 0 0 2
151 63
83 63
1 0 11 0 0 4096 0 2 0 0 15 2
84 114
132 114
2 1 11 0 0 8320 0 3 4 0 0 4
151 81
132 81
132 149
151 149
12
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 157
384 29 608 213
388 33 604 177
157 Inputs      Output
EN  D         Q
0   X    Q0 (no change)
1   0    0
1   1    1

"X" indicates "Don't care"
Q0 is state Q just prior
to EN going LOW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
460 179 492 203
464 183 488 199
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
190 178 222 202
194 182 218 198
3 (a)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
224 26 312 50
228 30 308 46
10 NAND LATCH
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
204 139 252 163
208 143 248 159
5 CLEAR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
204 125 252 149
208 129 248 145
5 _____
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
221 53 253 77
225 57 249 73
3 SET
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
221 39 253 63
225 43 249 59
3 ___
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
346 62 362 86
350 66 358 82
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
346 130 362 154
350 134 358 150
1 Q
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
346 122 362 146
350 126 358 142
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 63
196 243 420 307
200 247 416 295
63 D Latch (Transparent Latch)
  (a) structure
  (b) truth table
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 4.6e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
