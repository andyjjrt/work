CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 430
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 430
8912914 0
0
6 Title:
5 Name:
0
0
0
12
9 Terminal~
194 392 107 0 1 3
0 2
0
0 0 49504 270
8 OverTemp
6 -4 62 4
2 T1
-7 -25 7 -17
0
9 OverTemp;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
8953 0 0
0
0
2 +V
167 350 54 0 1 3
0 4
0
0 0 53600 0
3 +5V
-10 -14 11 -6
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
2 +V
167 287 55 0 1 3
0 6
0
0 0 53600 0
3 +5V
-11 -15 10 -7
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
7 Ground~
168 287 135 0 1 3
0 3
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 195 255 0 1 3
0 3
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
2 +V
167 112 93 0 1 3
0 8
0
0 0 53600 0
3 +5V
-10 -14 11 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
7 Ground~
168 133 200 0 1 3
0 3
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
12 Comparator5~
219 287 106 0 5 11
0 7 5 6 3 2
0
0 0 320 0
5 LM339
8 -16 43 -8
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP14
26

0 5 4 3 12 2 5 4 3 12
2 7 6 3 12 1 9 8 3 12
14 11 10 3 12 13 917522
88 0 0 0 4 1 1 0
1 U
3747 0 0
0
0
5 RRECT
94 133 157 0 2 5
0 7 3
5 RRECT
1 0 1088 0
2 1V
-7 -25 7 -17
2 U2
40 2 54 10
4 LM34
-13 3 15 11
0
28 %D %1 %2 DC 0 PWL( 0 0 10 2)
0
0
0
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
9 Resistor~
219 350 80 0 3 5
0 4 2 1
0
0 0 864 270
3 10k
7 0 28 8
2 Rp
11 -11 25 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 195 222 0 4 5
0 5 3 0 -1
0
0 0 864 270
2 2k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 195 165 0 3 5
0 8 5 1
0
0 0 864 270
2 8k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
12
1 0 2 0 0 4096 0 1 0 0 3 2
380 106
350 106
1 1 4 0 0 4224 0 2 10 0 0 2
350 63
350 62
5 2 2 0 0 4224 0 8 10 0 0 3
305 106
350 106
350 98
0 2 5 0 0 8320 0 0 8 11 0 4
195 193
251 193
251 100
269 100
1 3 6 0 0 4224 0 3 8 0 0 2
287 64
287 93
1 4 3 0 0 4224 0 4 8 0 0 2
287 129
287 119
1 1 7 0 0 8320 0 9 8 0 0 3
133 142
133 112
269 112
0 1 8 0 0 4224 0 0 12 9 0 3
112 131
195 131
195 147
1 0 8 0 0 0 0 6 0 0 0 2
112 102
112 148
1 2 3 0 0 0 0 5 11 0 0 2
195 249
195 240
2 1 5 0 0 0 0 12 11 0 0 2
195 183
195 204
1 2 3 0 0 0 0 7 9 0 0 2
133 194
133 186
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
128 92 184 112
132 96 181 110
7 10mV/�F
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 76
328 242 584 306
332 246 580 294
76 A temperature-limit detector 
using an LM339 analog voltage 
comparator.
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
267780172 8525888 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 1e-006 2
2
221 112
0 7 0 0 2	0 7 0 0
367 106
0 2 0 0 1	0 1 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 3 0 0
200 112
0 7 0 0 2	0 7 0 0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
