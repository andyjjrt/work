CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 458
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 458
8912914 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 125 88 0 1 11
0 11
0
0 0 21616 0
2 0V
-6 -16 8 -8
3 VIN
-36 -4 -15 4
1 A
-23 -5 -16 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 129 224 0 1 11
0 8
0
0 0 21616 0
2 0V
-6 -16 8 -8
4 VIN1
-39 -4 -11 4
1 B
-22 -5 -15 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
12 P-EMOS 3T:A~
219 323 97 0 3 7
0 7 8 9
0
0 0 1104 180
4 PMOS
18 0 46 8
2 Q1
18 -5 32 3
2 Q1
-36 -5 -22 3
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 2 3 1 2 3 1 0
109 0 0 0 0 0 0 0
1 Q
3618 0 0
0
0
12 P-EMOS 3T:A~
219 242 97 0 3 7
0 7 11 9
0
0 0 1104 692
4 PMOS
18 0 46 8
2 Q5
18 -5 32 3
2 Q1
18 -5 32 3
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 2 3 1 2 3 1 0
109 0 0 0 0 0 0 0
1 Q
6153 0 0
0
0
7 Ground~
168 280 261 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
2 +V
167 280 47 0 1 3
0 9
0
0 0 54384 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
4 +VDD
-12 -14 16 -6
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
12 N-EMOS 3T:A~
219 274 161 0 3 7
0 7 11 10
0
0 0 1104 0
4 NMOS
18 0 46 8
2 Q6
18 -5 32 3
2 Q2
18 -5 32 3
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 1 2 3 1 2 3 0
77 0 0 0 0 0 0 0
1 Q
9914 0 0
0
0
12 N-EMOS 3T:A~
219 274 215 0 3 7
0 10 8 2
0
0 0 1104 0
4 NMOS
18 0 46 8
2 Q2
18 -5 32 3
2 Q2
18 -5 32 3
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 1 2 3 1 2 3 0
77 0 0 0 0 0 0 0
1 Q
3747 0 0
0
0
11 Multimeter~
205 446 110 0 21 21
0 7 12 13 2 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
7 Ground~
168 471 148 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7931 0 0
0
0
17
0 0 1 0 0 4272 0 0 0 4 3 2
505 204
505 283
0 0 3 0 0 4240 0 0 0 0 0 2
461 208
461 279
0 0 4 0 0 4240 0 0 0 0 0 2
424 283
547 283
0 0 5 0 0 4240 0 0 0 0 0 2
423 204
546 204
0 0 6 0 0 4240 0 0 0 0 0 2
423 219
546 219
1 4 2 0 0 4096 0 10 9 0 0 2
471 142
471 133
0 1 7 0 0 4224 0 0 9 11 0 2
280 133
421 133
0 2 8 0 0 12416 0 0 3 15 0 5
205 224
205 281
350 281
350 88
337 88
1 0 9 0 0 4096 0 6 0 0 10 2
280 56
280 71
3 3 9 0 0 8320 0 4 3 0 0 4
248 79
248 71
313 71
313 79
1 0 7 0 0 0 0 7 0 0 12 2
280 143
280 123
1 1 7 0 0 0 0 4 3 0 0 4
248 115
248 123
313 123
313 115
3 1 2 0 0 4224 0 8 5 0 0 2
280 233
280 255
3 1 10 0 0 4224 0 7 8 0 0 2
280 179
280 197
2 1 8 0 0 0 0 8 2 0 0 2
256 224
141 224
0 2 11 0 0 4096 0 0 7 17 0 3
205 88
205 170
256 170
1 2 11 0 0 4224 0 1 4 0 0 2
137 88
224 88
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 81
421 200 557 304
425 204 553 284
81  A    B     X
LOW  LOW   HIGH
LOW  HIGH  HIGH
HIGH LOW   HIGH
HIGH HIGH  HIGH
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
221 307 349 331
225 311 345 327
15 CMOS NAND gate.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
375 99 399 123
379 103 395 119
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
359 113 399 137
363 117 395 133
4 X=AB
0
1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
-1241054938 1210432 100 100 0 0
77 66 587 246
420 103 581 173
587 66
77 66
587 66
587 246
0 0
0.003 0 5.4 0 0.003 5.4
12401 0
4 1e-007 2
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
