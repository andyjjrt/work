CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 440
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 440
11010066 0
0
6 Title:
5 Name:
0
0
0
5
9 Terminal~
194 365 157 0 1 3
0 2
0
0 0 49520 270
4 Vout
7 -4 35 4
2 T1
-7 -25 7 -17
0
5 Vout;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
8953 0 0
0
0
7 Ground~
168 220 231 0 1 3
0 3
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4441 0 0
0
0
10 Capacitor~
219 220 200 0 2 5
0 4 3
0
0 0 848 270
3 1uF
11 0 32 8
1 C
18 -10 25 -2
0
0
18 %D %1 %2 %V IC=.8V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3618 0 0
0
0
5 7414~
219 271 156 0 2 22
0 4 2
0
0 0 368 0
6 74LS14
1 9 43 17
3 U1A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 1 0
1 U
6153 0 0
0
0
9 Resistor~
219 220 121 0 2 5
0 2 4
0
0 0 880 270
4 1.2k
8 0 36 8
1 R
18 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
5
1 0 2 0 0 4096 0 1 0 0 3 2
353 156
321 156
1 0 4 0 0 4096 0 4 0 0 5 2
256 156
220 156
1 2 2 0 0 8336 0 5 4 0 0 5
220 103
220 92
321 92
321 156
292 156
2 1 3 0 0 4224 0 3 2 0 0 2
220 209
220 225
2 1 4 0 0 4224 0 5 3 0 0 2
220 139
220 191
1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 98
103 279 511 323
107 283 507 315
98 Schmitt-trigger oscillator using a 7414 INVERTER. 
A 7413 Schmitt-trigger NAND may also be used.
0
16 2 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.006 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1434845562 8550464 100 100 0 0
77 66 587 156
4 440 635 663
422 66
306 66
587 66
587 156
0 0
0.00405882 0.00269412 4.2 0 0.006 0.006
12401 0
4 0.001 2
2
339 156
0 2 0 0 1	0 1 0 0
239 156
0 4 0 0 1	0 2 0 0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
