CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 393
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 393 635 502
25165842 0
0
6 Title:
5 Name:
0
0
0
5
5 SCOPE
12 158 74 0 1 11
0 3
0
0 0 57584 0
1 A
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SCOPE
12 193 74 0 1 11
0 2
0
0 0 57584 0
1 B
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 291 74 0 1 11
0 4
0
0 0 57584 0
3 Out
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 4001~
219 225 129 0 3 22
0 3 2 4
0
0 0 112 0
4 4001
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
6153 0 0
0
0
9 Data Seq~
170 97 84 0 17 18
0 9 10 11 12 13 14 2 3 15
16 17 1 20 10 1 0 33
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
5394 0 0
0
0
AAACACADABAAACADABAAACACACACACACACACACACACACACACACACACACACACACACAC
10
1 0 2 0 0 4112 0 2 0 0 4 2
193 86
193 138
1 0 3 0 0 4112 0 1 0 0 3 2
158 86
158 120
1 8 3 0 0 4240 0 4 5 0 0 2
212 120
129 120
2 7 2 0 0 4240 0 4 5 0 0 4
212 138
144 138
144 111
129 111
3 1 4 0 0 8336 0 4 3 0 0 3
264 129
291 129
291 86
0 0 5 0 0 4224 0 0 0 0 0 5
303 223
572 223
572 256
303 256
303 223
0 0 1 0 0 4256 0 0 0 0 0 2
450 58
450 144
0 0 6 0 0 4224 0 0 0 0 0 2
394 144
486 144
0 0 7 0 0 4224 0 0 0 0 0 2
394 77
486 77
0 0 8 0 0 4224 0 0 0 0 0 2
394 58
486 58
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
254 140 302 164
258 144 298 160
5 x=A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
271 125 303 149
275 129 299 145
3 ___
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
305 220 571 257
309 224 568 252
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
44 228 252 252
48 232 248 248
25 NOR gate and truth table.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 59
391 58 487 162
395 62 483 142
59 A   B   A+B
0   0    1
0   1    0
1   0    0
1   1    0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
455 44 487 68
459 48 483 64
3 ___
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 2e-005 1e-008 1e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
