CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 458
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 458
8912914 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 76 193 0 1 11
0 4
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
3 VIN
-39 -3 -18 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
9 Terminal~
194 176 160 0 1 3
0 2
0
0 0 49520 270
4 VOUT
-8 6 20 14
2 T1
-7 -25 7 -17
0
5 VOUT;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
1 T
4441 0 0
0
0
10 N-EMOS 3T~
219 120 184 0 3 7
0 2 4 3
0
0 0 80 0
6 2N3797
10 -4 52 4
2 Q1
23 -14 37 -6
0
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 2 3 1 2 3 1 0
77 0 0 0 1 0 0 0
1 Q
3618 0 0
0
0
10 N-EMOS 3T~
219 120 133 0 3 7
0 5 5 2
0
0 0 80 0
4 NMOS
17 -4 45 4
2 Q6
23 -14 37 -6
0
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 1 2 3 1 2 3 0
77 0 0 0 1 0 0 0
1 Q
6153 0 0
0
0
2 +V
167 126 80 0 1 3
0 5
0
0 0 54128 0
3 +5V
6 -3 27 5
3 VDD
-9 -15 12 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
7 Ground~
168 126 217 0 1 3
0 3
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 214 182 0 1 3
0 3
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
11 Multimeter~
205 189 130 0 21 21
0 2 12 13 3 0 0 0 0 0
32 52 46 57 51 48 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
15
1 0 2 0 0 0 0 2 0 0 4 2
164 159
164 159
2 1 4 0 0 4224 0 3 1 0 0 2
102 193
88 193
2 0 5 0 0 8320 0 4 0 0 7 4
102 142
90 142
90 102
126 102
1 0 2 0 0 8320 0 8 0 0 6 3
164 153
164 159
126 159
1 4 3 0 0 4224 0 7 8 0 0 2
214 176
214 153
3 1 2 0 0 0 0 4 3 0 0 2
126 151
126 166
1 1 5 0 0 0 0 5 4 0 0 2
126 89
126 115
1 3 3 0 0 0 0 6 3 0 0 2
126 211
126 202
0 0 6 0 0 4224 0 0 0 0 0 2
471 127
471 190
0 0 7 0 0 4224 0 0 0 0 0 2
417 127
417 190
0 0 1 0 0 4256 0 0 0 0 0 2
367 124
367 194
0 0 8 0 0 4224 0 0 0 0 0 2
299 194
554 194
0 0 9 0 0 4224 0 0 0 0 0 2
298 166
553 166
0 0 10 0 0 4224 0 0 0 0 0 2
297 124
552 124
0 0 11 0 0 4224 0 0 0 0 0 2
297 138
552 138
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
210 293 330 317
214 297 326 313
14 N-MOS INVERTER
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 178
295 119 554 207
299 123 551 193
178    VIN      Q1      Q2    VOUT = VIN
0V         RON =  ROFF =    +5V
(logic 0)  100k    10     (logic 1)
+5V        RON =  RON =    +0.05V
(logic 1)  100k    1k     (logic 0)
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
441 144 462 164
445 148 459 162
2 10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
404 234 436 258
408 238 432 254
3 (b)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
108 234 140 258
112 238 136 254
3 (a)
0
1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1605960484 1210432 100 100 0 0
77 66 587 246
346 102 507 172
587 66
77 66
587 66
587 246
0 0
0.003 0 5.4 0 0.003 5.4
12401 0
4 2 2
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
