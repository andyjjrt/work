CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 436 635 675
27262994 0
0
6 Title:
5 Name:
0
0
0
13
5 SCOPE
12 162 110 0 1 11
0 11
0
0 0 57584 0
2 CP
-8 -4 6 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SCOPE
12 456 62 0 1 11
0 3
0
0 0 57584 0
2 Q0
-8 -4 6 4
3 U11
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 436 47 0 1 11
0 4
0
0 0 57584 0
2 Q1
-8 -4 6 4
3 U10
-11 -14 10 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 417 62 0 1 11
0 5
0
0 0 57584 0
2 Q2
-8 -4 6 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
5 SCOPE
12 397 47 0 1 11
0 6
0
0 0 57584 0
2 Q3
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 377 62 0 1 11
0 7
0
0 0 57584 0
2 Q4
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 358 47 0 1 11
0 8
0
0 0 57584 0
2 Q5
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 339 62 0 1 11
0 9
0
0 0 57584 0
2 Q6
-8 -4 6 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 319 47 0 1 11
0 10
0
0 0 57584 0
2 Q7
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
7 Pulser~
4 106 130 0 10 12
0 14 15 11 16 0 0 5 5 6
7
0
0 0 4144 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7931 0 0
0
0
2 +V
167 215 72 0 1 3
0 12
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
9 Inverter~
13 190 139 0 2 22
0 10 13
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8903 0 0
0
0
7 74LS164
127 259 121 0 12 25
0 12 12 11 13 10 9 8 7 6
5 4 3
0
0 0 4464 0
8 74ALS164
-28 -51 28 -43
2 U1
-7 -52 7 -44
0
15 DVCC=14;DGND=7;
96 %D [%14bi %7bi %1i %2i %3i %4i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o] %M
0
12 type:digital
5 DIP14
25

0 1 2 8 9 13 12 11 10 6
5 4 3 1 2 8 9 13 12 11
10 6 5 4 3 0
65 0 0 0 1 0 0 0
1 U
3834 0 0
0
0
15
0 0 2 0 0 4224 0 0 0 0 0 5
305 268
576 268
576 301
305 301
305 268
12 1 3 0 0 4224 0 13 2 0 0 3
291 157
456 157
456 74
11 1 4 0 0 4224 0 13 3 0 0 3
291 148
436 148
436 59
10 1 5 0 0 4224 0 13 4 0 0 3
291 139
417 139
417 74
9 1 6 0 0 4224 0 13 5 0 0 3
291 130
397 130
397 59
8 1 7 0 0 4224 0 13 6 0 0 3
291 121
377 121
377 74
7 1 8 0 0 4224 0 13 7 0 0 3
291 112
358 112
358 59
6 1 9 0 0 4224 0 13 8 0 0 3
291 103
339 103
339 74
5 1 10 0 0 8192 0 13 9 0 0 3
291 94
319 94
319 59
1 0 11 0 0 4096 0 1 0 0 11 2
162 122
162 121
3 3 11 0 0 4224 0 10 13 0 0 2
130 121
227 121
1 0 12 0 0 4096 0 13 0 0 13 2
227 94
215 94
1 2 12 0 0 4224 0 11 13 0 0 3
215 81
215 103
227 103
0 1 10 0 0 8320 0 0 12 9 0 5
303 94
303 174
162 174
162 139
175 139
2 4 13 0 0 4224 0 12 13 0 0 2
211 139
221 139
2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 63
26 251 226 315
30 255 222 303
63 The 74ALS164 8-bit 
serial in/parallel out 
shift register.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
307 265 573 302
311 269 570 297
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 2
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.003 2e-006 2e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
619643552 1210432 100 100 0 0
77 66 587 156
11 95 172 165
587 66
77 66
587 66
587 156
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 1 0.001
0
387777332 8550464 100 100 0 0
77 66 587 246
3 436 635 771
442 66
170 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
13425 0
2 0.0005 5
3
323 159
0 5 0 59 2	0 2 0 0
331 150
0 4 0 30 1	0 16 0 0
337 141
0 3 0 0 1	0 3 0 0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
