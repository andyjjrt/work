CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 420
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 420
8388626 0
0
6 Title:
5 Name:
0
0
0
7
13 Logic Switch~
5 82 142 0 1 11
0 10
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
5 Clock
-56 -3 -21 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 131 189 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21600 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
5 Reset
-52 -5 -17 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 131 158 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21600 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 K
-26 -4 -19 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 131 126 0 1 11
0 8
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 J
-26 -4 -19 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 131 95 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21600 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
3 Set
-39 -4 -18 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5394 0 0
0
0
14 Logic Display~
6 259 111 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
6 74112~
219 198 169 0 7 32
0 9 8 10 7 6 11 5
0
0 0 4192 0
7 74LS112
-3 -60 46 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 1 0
1 U
9914 0 0
0
0
10
0 0 2 0 0 4224 0 0 0 0 0 2
311 95
560 95
0 0 1 0 0 4256 0 0 0 1 0 2
400 95
400 176
0 0 3 0 0 4224 0 0 0 0 0 2
311 176
560 176
0 0 4 0 0 4224 0 0 0 0 0 2
311 111
560 111
1 7 5 0 0 8320 0 6 7 0 0 3
259 129
259 133
222 133
1 5 6 0 0 4224 0 2 7 0 0 3
143 189
198 189
198 181
1 4 7 0 0 4224 0 3 7 0 0 4
143 158
160 158
160 151
174 151
1 2 8 0 0 4224 0 4 7 0 0 4
143 126
160 126
160 133
174 133
1 1 9 0 0 4224 0 5 7 0 0 3
143 95
198 95
198 106
3 1 10 0 0 4224 0 7 1 0 0 2
168 142
94 142
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 47
100 264 484 288
104 268 480 284
47 Clocked J-K flip-flop with asynchronous inputs.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 156
301 92 573 216
305 96 569 192
156  SET  RESET    FF response
  1     1    Clocked operation*
  0     1    Q = 1
  1     0    Q = 0
  1     1    Not used
 *Q will respond to J, K, and CP
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
309 79 341 103
313 83 337 99
3 ___
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
349 79 397 103
353 83 393 99
5 _____
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
88 72 116 92
92 76 113 90
3 ___
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
76 165 118 185
80 169 115 183
5 _____
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 3.2e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
0.016 0 24 0 0.016 24
12401 0
0 2 2
0
0 0 100 100 0 0
77 66 587 246
0 0 0 0
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547059 4.8 1.70667 0.003 0.003
12401 0
0 0.001 2
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
