CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 21 100 9
4 70 635 393
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 393
8388626 0
0
6 Title:
5 Name:
0
0
0
6
5 4049~
219 201 159 0 2 22
0 5 3
0
0 0 96 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 1 3 0
1 U
8953 0 0
0
0
14 Logic Display~
6 326 93 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
5 4023~
219 273 120 0 4 22
0 6 4 3 2
0
0 0 96 0
4 4023
-14 -28 14 -20
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
3618 0 0
0
0
13 Logic Switch~
5 149 159 0 1 11
0 5
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 C
-24 -3 -17 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 149 129 0 1 11
0 4
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 B
-23 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 149 103 0 1 11
0 6
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-24 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7734 0 0
0
0
5
1 4 2 0 0 16 0 2 3 0 0 3
326 111
326 120
300 120
3 2 3 0 0 16 0 3 1 0 0 4
249 129
240 129
240 159
222 159
2 1 4 0 0 16 0 3 5 0 0 4
249 120
201 120
201 129
161 129
1 1 5 0 0 16 0 1 4 0 0 2
186 159
161 159
1 1 6 0 0 16 0 3 6 0 0 4
249 111
201 111
201 103
161 103
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
210 242 378 266
214 246 374 262
20 DeMorgan's theorems.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
224 139 240 163
228 143 236 159
1 C
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
224 131 240 155
228 135 236 151
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
448 127 464 151
452 131 460 147
1 _
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
480 129 512 153
484 133 508 149
3 _ _
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
416 129 464 153
420 133 460 149
5 _ _ _
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
385 129 401 153
389 133 397 149
1 _
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
353 127 401 151
357 131 397 147
5 _____
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 25
320 143 528 167
324 147 524 163
25 z = A�B�C = A+B+C = A+B+C
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 2e-005 1e-008 1e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
