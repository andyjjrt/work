CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 440
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 440 635 612
27262994 0
0
6 Title:
5 Name:
0
0
0
22
13 Logic Switch~
5 130 116 0 1 11
0 6
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
7 DATA IN
-66 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
14 Logic Display~
6 538 43 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 465 43 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 387 43 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 309 43 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 234 43 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
5 SCOPE
12 182 161 0 1 11
0 8
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 211 49 0 1 11
0 6
0
0 0 57568 0
3 DIN
-11 -4 10 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
5 SCOPE
12 286 49 0 1 11
0 5
0
0 0 57568 0
2 X3
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
5 SCOPE
12 364 49 0 1 11
0 4
0
0 0 57568 0
2 X2
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7931 0 0
0
0
5 SCOPE
12 442 49 0 1 11
0 3
0
0 0 57568 0
2 X1
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9325 0 0
0
0
5 SCOPE
12 515 49 0 1 11
0 2
0
0 0 57568 0
2 X0
-8 -4 6 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8903 0 0
0
0
2 +V
167 480 81 0 1 3
0 9
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3834 0 0
0
0
2 +V
167 402 82 0 1 3
0 10
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
2 +V
167 325 82 0 1 3
0 11
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7668 0 0
0
0
2 +V
167 247 81 0 1 3
0 12
0
0 0 53472 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
6 74113~
219 480 133 0 6 22
0 3 8 13 9 17 2
0
0 0 4192 0
7 74LS113
-25 -42 24 -34
3 U2B
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 512 2 2 2 0
1 U
3874 0 0
0
0
6 74113~
219 402 133 0 6 22
0 4 8 14 10 13 3
0
0 0 4192 0
7 74LS113
-25 -42 24 -34
3 U2A
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 1 2 0
1 U
6671 0 0
0
0
6 74113~
219 325 133 0 6 22
0 5 8 15 11 14 4
0
0 0 4192 0
7 74LS113
-25 -42 24 -34
3 U1B
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 11 13 12 10 8 9 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 2 1 0
1 U
3789 0 0
0
0
6 74113~
219 247 133 0 6 22
0 6 8 16 12 15 5
0
0 0 4192 0
7 74LS113
-25 -42 24 -34
3 U1A
-11 24 10 32
0
15 DVCC=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
19

0 3 1 2 4 6 5 3 1 2
4 6 5 11 13 12 10 8 9 0
65 0 0 0 2 1 1 0
1 U
4871 0 0
0
0
9 Inverter~
13 183 134 0 2 22
0 6 16
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3750 0 0
0
0
7 Pulser~
4 125 183 0 10 12
0 18 19 8 20 0 0 5 5 6
7
0
0 0 4128 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8778 0 0
0
0
29
0 0 7 0 0 16 0 0 0 0 0 5
307 279
578 279
578 310
307 310
307 279
1 0 2 0 0 4096 0 2 0 0 7 2
538 61
515 61
1 0 3 0 0 4096 0 3 0 0 8 2
465 61
442 61
1 0 4 0 0 4096 0 4 0 0 9 2
387 61
364 61
1 0 5 0 0 4096 0 5 0 0 10 2
309 61
286 61
1 0 6 0 0 4096 0 6 0 0 11 2
234 61
211 61
1 6 2 0 0 4224 0 12 17 0 0 3
515 61
515 116
504 116
1 0 3 0 0 4224 0 11 0 0 23 2
442 61
442 116
1 0 4 0 0 4224 0 10 0 0 25 2
364 61
364 116
1 0 5 0 0 4224 0 9 0 0 27 2
286 61
286 116
1 0 6 0 0 4096 0 8 0 0 28 2
211 61
211 116
1 0 8 0 0 4096 0 7 0 0 21 2
182 173
182 174
1 4 9 0 0 4224 0 13 17 0 0 2
480 90
480 89
1 4 10 0 0 4224 0 14 18 0 0 2
402 91
402 89
1 4 11 0 0 4224 0 15 19 0 0 2
325 91
325 89
1 4 12 0 0 4224 0 16 20 0 0 2
247 90
247 89
1 0 6 0 0 0 0 21 0 0 28 3
168 134
152 134
152 116
2 0 8 0 0 8192 0 20 0 0 21 3
216 125
211 125
211 174
2 0 8 0 0 0 0 19 0 0 21 3
294 125
286 125
286 174
2 0 8 0 0 0 0 18 0 0 21 3
371 125
364 125
364 174
3 2 8 0 0 4224 0 22 17 0 0 4
149 174
443 174
443 125
449 125
5 3 13 0 0 4224 0 18 17 0 0 2
432 134
456 134
6 1 3 0 0 0 0 18 17 0 0 2
426 116
456 116
5 3 14 0 0 4224 0 19 18 0 0 2
355 134
378 134
6 1 4 0 0 0 0 19 18 0 0 2
349 116
378 116
5 3 15 0 0 4224 0 20 19 0 0 2
277 134
301 134
6 1 5 0 0 0 0 20 19 0 0 2
271 116
301 116
1 1 6 0 0 4224 0 1 20 0 0 2
142 116
223 116
2 3 16 0 0 4224 0 21 20 0 0 2
204 134
223 134
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
309 276 575 313
313 280 572 308
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 4
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 24
46 283 246 307
50 287 242 303
24 Four-bit shift register.
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
