CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 436 635 590
27262994 0
0
6 Title:
5 Name:
0
0
0
11
7 Pulser~
4 67 178 0 10 12
0 10 11 8 12 0 0 20 20 19
7
0
0 0 1056 0
0
2 V1
-7 -28 7 -20
5 Clock
-17 -28 18 -20
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 1 0 0
1 V
8953 0 0
0
0
14 Logic Display~
6 395 69 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 311 69 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 228 69 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
5 SCOPE
12 115 149 0 1 11
0 8
0
0 0 57568 0
2 CP
-8 -4 6 4
2 U9
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
5 SCOPE
12 205 75 0 1 11
0 7
0
0 0 57568 0
2 Q2
-8 -4 6 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
5 SCOPE
12 288 75 0 1 11
0 6
0
0 0 57568 0
2 Q1
-8 -4 6 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
5 SCOPE
12 372 75 0 1 11
0 5
0
0 0 57568 0
2 Q0
-8 -4 6 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3747 0 0
0
0
12 D Flip-Flop~
219 338 161 0 4 9
0 6 8 9 5
0
0 0 4192 0
3 DFF
-10 -53 11 -45
2 U3
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3549 0 0
0
0
12 D Flip-Flop~
219 254 161 0 4 9
0 7 8 13 6
0
0 0 4192 0
3 DFF
-10 -53 11 -45
2 U2
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
12 D Flip-Flop~
219 171 161 0 4 9
0 9 8 14 7
0
0 0 4192 0
3 DFF
-10 -53 11 -45
2 U1
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9325 0 0
0
0
18
0 0 2 0 0 16 0 0 0 0 0 5
315 276
586 276
586 308
315 308
315 276
0 0 1 0 0 4256 0 0 0 4 3 2
508 18
508 243
0 0 2 0 0 4224 0 0 0 0 0 2
442 243
552 243
0 0 3 0 0 4224 0 0 0 0 0 2
442 18
552 18
0 0 4 0 0 4224 0 0 0 0 0 2
441 50
551 50
1 0 5 0 0 4096 0 2 0 0 16 2
395 87
372 87
1 0 6 0 0 4096 0 3 0 0 9 2
311 87
288 87
1 0 7 0 0 4096 0 4 0 0 10 2
228 87
205 87
1 0 6 0 0 4224 0 7 0 0 17 2
288 87
288 125
1 0 7 0 0 4224 0 6 0 0 18 2
205 87
205 125
1 0 8 0 0 4096 0 5 0 0 15 2
115 161
115 169
3 1 9 0 0 12416 0 9 11 0 0 6
368 143
385 143
385 102
139 102
139 125
147 125
2 0 8 0 0 8192 0 11 0 0 15 3
147 143
136 143
136 169
2 0 8 0 0 0 0 10 0 0 15 3
230 143
223 143
223 169
3 2 8 0 0 4224 0 1 9 0 0 4
91 169
308 169
308 143
314 143
4 1 5 0 0 8320 0 9 8 0 0 3
362 125
372 125
372 87
4 1 6 0 0 0 0 10 9 0 0 2
278 125
314 125
4 1 7 0 0 0 0 11 10 0 0 2
195 125
230 125
3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
317 273 583 310
321 277 580 305
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 22
61 281 245 305
65 285 241 301
22 Four-bit ring counter.
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 198
436 14 564 298
440 18 560 242
198          CLOCK
Q2 Q1 Q0 pulse
0  0  0    0
1  0  0    1
1  1  0    2
1  1  1    3
0  1  1    4
0  0  1    5
0  0  0    6
1  0  0    7
1  1  0    8
.  .  .    .
.  .  .    .
.  .  .    .
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.003 6e-006 6e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
62522106 8550464 100 100 0 0
77 66 587 246
3 436 635 771
451 66
213 66
587 66
587 246
0 0
0.0022 0.0008 30 -30 0.003 0.003
13425 0
2 0.0005 10
5
182 159
0 8 0 60 1	0 18 0 0
385 141
0 5 0 -59 1	0 15 0 0
375 150
0 4 0 -29 1	0 19 0 0
363 159
0 3 0 0 1	0 17 0 0
352 168
0 2 0 32 1	0 19 0 0
110889084 8550464 100 100 0 0
77 66 587 246
3 436 635 771
442 66
170 66
587 66
587 182
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2
1
348 141
0 4 0 0 1	0 17 0 0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
