CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 742
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 742
8912914 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 177 446 0 1 11
0 4
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
11 Input A (1)
-97 -3 -20 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 155 185 0 1 11
0 9
0
0 0 21600 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
11 Input A (1)
-96 -3 -19 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
11 Multimeter~
205 449 421 0 21 21
0 3 16 17 2 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 82
0
0 0 16448 0
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
3618 0 0
0
0
7 Ground~
168 474 462 0 1 3
0 2
0
0 0 53344 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
6 Diode~
219 219 469 0 2 5
0 2 4
0
0 0 64 90
5 DIODE
11 0 46 8
2 D4
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
5394 0 0
0
0
6 Diode~
219 219 424 0 2 5
0 4 5
0
0 0 64 90
5 DIODE
11 0 46 8
2 D3
22 -10 36 -2
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7734 0 0
0
0
7 Ground~
168 294 505 0 1 3
0 2
0
0 0 54368 0
0
4 GND3
-14 -26 14 -18
7 GND (7)
12 -1 61 7
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9914 0 0
0
0
2 +V
167 294 384 0 1 3
0 5
0
0 0 54368 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
9 +VDD (14)
7 -3 70 5
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3747 0 0
0
0
12 P-EMOS 3T:A~
219 288 421 0 3 7
0 3 4 5
0
0 0 1088 692
4 PMOS
18 0 46 8
2 Q5
18 -5 32 3
2 Q1
18 -5 32 3
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
109 0 0 0 1 0 0 0
1 Q
3549 0 0
0
0
12 N-EMOS 3T:A~
219 288 473 0 3 7
0 3 4 2
0
0 0 1088 0
4 NMOS
18 0 46 8
2 Q6
18 -5 32 3
2 Q2
18 -5 32 3
0
17 %D %1 %2 %3 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
77 0 0 0 1 0 0 0
1 Q
7931 0 0
0
0
7 Ground~
168 496 217 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9325 0 0
0
0
11 Multimeter~
205 471 176 0 21 21
0 7 18 19 2 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 82
0
0 0 16448 0
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
7 Ground~
168 290 297 0 1 3
0 2
0
0 0 54368 0
0
4 GND1
-14 -26 14 -18
7 GND (7)
12 -1 61 7
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3834 0 0
0
0
2 +V
167 147 87 0 1 3
0 8
0
0 0 54368 90
2 5V
-7 -15 7 -7
2 V1
-7 -25 7 -17
9 +Vcc (14)
-73 -6 -10 2
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
6 Diode~
219 185 256 0 2 5
0 2 9
0
0 0 576 90
5 DIODE
11 0 46 8
2 D1
12 -5 26 3
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
7668 0 0
0
0
12 NPN Trans:B~
219 311 228 0 3 7
0 7 10 2
0
0 0 576 0
3 NPN
17 0 38 8
2 Q3
8 -3 22 5
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
4718 0 0
0
0
6 Diode~
219 316 184 0 2 5
0 13 7
0
0 0 576 270
5 DIODE
11 0 46 8
2 D2
12 -5 26 3
0
0
11 %D %1 %2 %M
0
0
8 DIODE0.4
5

0 -54 -44 -54 -44 0
68 0 0 0 1 0 0 0
1 D
3874 0 0
0
0
12 NPN Trans:B~
219 311 152 0 3 7
0 14 11 13
0
0 0 576 0
3 NPN
17 0 38 8
2 Q4
9 -2 23 6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
6671 0 0
0
0
12 NPN Trans:B~
219 259 185 0 3 7
0 11 12 10
0
0 0 576 0
3 NPN
17 0 38 8
2 Q2
8 -1 22 7
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
3789 0 0
0
0
12 NPN Trans:B~
219 218 178 0 3 7
0 12 15 9
0
0 0 576 270
3 NPN
-13 30 8 38
2 Q1
-9 12 5 20
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 0
81 0 0 0 1 1 0 0
1 Q
4871 0 0
0
0
9 Resistor~
219 264 257 0 4 5
0 10 2 0 -1
0
0 0 864 270
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3750 0 0
0
0
9 Resistor~
219 316 110 0 3 5
0 8 14 1
0
0 0 864 270
3 115
7 0 28 8
2 R4
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8778 0 0
0
0
9 Resistor~
219 264 111 0 3 5
0 8 11 1
0
0 0 864 270
4 1.6k
8 0 36 8
2 R2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
538 0 0
0
0
9 Resistor~
219 216 114 0 3 5
0 8 15 1
0
0 0 864 270
4 3.6k
8 0 36 8
2 R1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6843 0 0
0
0
31
1 0 3 0 0 8320 0 3 0 0 9 3
424 444
424 447
294 447
1 4 2 0 0 4096 0 4 3 0 0 2
474 456
474 444
1 0 4 0 0 4096 0 6 0 0 5 2
219 434
219 446
2 0 4 0 0 4096 0 5 0 0 5 2
219 459
219 446
1 0 4 0 0 4224 0 1 0 0 8 2
189 446
262 446
1 0 2 0 0 8192 0 5 0 0 11 3
219 479
219 494
294 494
2 0 5 0 0 8320 0 6 0 0 10 3
219 414
219 399
294 399
2 2 4 0 0 0 0 9 10 0 0 4
270 412
262 412
262 482
270 482
1 1 3 0 0 0 0 9 10 0 0 2
294 439
294 455
1 3 5 0 0 0 0 8 9 0 0 2
294 393
294 403
1 3 2 0 0 0 0 7 10 0 0 2
294 499
294 491
0 0 6 0 0 4224 0 0 0 0 0 3
124 198
124 227
117 227
1 0 7 0 0 8320 0 12 0 0 27 3
446 199
446 202
316 202
1 4 2 0 0 0 0 11 12 0 0 2
496 211
496 199
1 0 8 0 0 4096 0 24 0 0 17 2
216 96
216 85
1 0 8 0 0 0 0 23 0 0 17 2
264 93
264 85
1 1 8 0 0 4224 0 14 22 0 0 3
158 85
316 85
316 92
2 0 9 0 0 4224 0 15 0 0 25 2
185 246
185 185
1 0 2 0 0 0 0 13 0 0 21 2
290 291
290 283
2 0 2 0 0 0 0 21 0 0 21 2
264 275
264 283
3 1 2 0 0 8320 0 16 15 0 0 4
316 246
316 283
185 283
185 266
2 0 10 0 0 4096 0 16 0 0 26 2
293 228
264 228
2 0 11 0 0 4096 0 18 0 0 30 2
293 152
264 152
1 2 12 0 0 4224 0 20 19 0 0 2
234 185
241 185
3 1 9 0 0 0 0 20 2 0 0 2
198 185
167 185
3 1 10 0 0 4224 0 19 21 0 0 2
264 203
264 239
2 1 7 0 0 0 0 17 16 0 0 2
316 194
316 210
3 1 13 0 0 4224 0 18 17 0 0 2
316 170
316 174
2 1 14 0 0 4224 0 22 18 0 0 2
316 128
316 134
2 1 11 0 0 4224 0 23 19 0 0 2
264 129
264 167
2 2 15 0 0 4224 0 24 20 0 0 2
216 132
216 162
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 91
67 575 491 619
71 579 487 611
91 (a) TTL INVERTER circuit; (b) CMOS INVERTER circuit.
Pin numbers are given in parentheses.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
343 184 434 204
347 188 431 202
12 Output Y (2)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
263 310 295 334
267 314 291 330
3 (a)
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
42 215 119 235
46 219 116 233
10 Pin number
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
117 189 133 213
121 193 129 209
1 ^
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
267 522 299 546
271 526 295 542
3 (b)
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
321 427 412 447
325 431 409 445
12 Output Y (2)
0
1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
928973094 1210432 100 100 0 0
0 0 0 0
8 92 169 162
0 0
0 0
0 0
0 0
0 0
0.016 0 24 0 0.016 24
12401 0
4 2 2
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 0.001 2e+012
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
