CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 436
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 436
10485778 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 85 218 0 1 11
0 4
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
3 MR1
-35 -5 -14 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 85 236 0 1 11
0 5
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
3 MR2
-36 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
7 Pulser~
4 56 154 0 10 12
0 14 15 16 3 0 0 20 20 21
7
0
0 0 560 0
0
3 CP0
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 1 0 0
1 V
3618 0 0
0
0
12 Hex Display~
7 541 49 0 16 19
10 2 8 7 6 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53360 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6153 0 0
0
0
6 74112~
219 184 181 0 7 32
0 13 13 3 13 9 17 2
0
0 0 4208 0
7 74LS112
-3 -60 46 -52
3 U2B
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 2 5 0
1 U
5394 0 0
0
0
14 Logic Display~
6 484 56 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 389 56 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
14 Logic Display~
6 300 58 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 214 58 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Q0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3549 0 0
0
0
2 +V
167 150 106 0 1 3
0 13
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7931 0 0
0
0
10 2-In NAND~
219 133 227 0 3 22
0 4 5 9
0
0 0 112 0
6 74LS00
-14 -24 28 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
9325 0 0
0
0
2 +V
167 234 107 0 1 3
0 12
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8903 0 0
0
0
6 74112~
219 268 182 0 7 32
0 12 12 2 12 9 18 8
0
0 0 4208 0
7 74LS112
-3 -60 46 -52
3 U1A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 7 0
1 U
3834 0 0
0
0
2 +V
167 323 108 0 1 3
0 11
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3363 0 0
0
0
6 74112~
219 357 183 0 7 32
0 11 11 8 11 9 19 7
0
0 0 4208 0
7 74LS112
-3 -60 46 -52
3 U1B
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 2 7 0
1 U
7668 0 0
0
0
2 +V
167 411 108 0 1 3
0 10
0
0 0 53488 0
2 5V
-7 -22 7 -14
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4718 0 0
0
0
6 74112~
219 445 183 0 7 32
0 10 10 7 10 9 20 6
0
0 0 4208 0
7 74LS112
-3 -60 46 -52
3 U3A
21 -61 42 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 8 0
1 U
3874 0 0
0
0
9 Terminal~
194 73 202 0 1 3
0 2
0
0 0 49520 90
3 CP1
-25 -6 -4 2
2 T1
-8 -25 6 -17
0
4 CP1;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
1 T
6671 0 0
0
0
31
3 4 3 0 0 4224 0 5 3 0 0 2
154 154
86 154
0 0 2 0 0 8192 0 0 0 5 19 3
104 200
104 92
214 92
1 1 4 0 0 4224 0 1 11 0 0 2
97 218
109 218
1 2 5 0 0 4224 0 2 11 0 0 2
97 236
109 236
1 3 2 0 0 4112 0 18 13 0 0 4
84 200
224 200
224 155
238 155
4 0 6 0 0 8192 0 4 0 0 10 3
532 73
532 77
484 77
3 0 7 0 0 8320 0 4 0 0 11 3
538 73
538 82
389 82
2 0 8 0 0 8320 0 4 0 0 12 3
544 73
544 87
300 87
1 0 2 0 0 8320 0 4 0 0 19 3
550 73
550 92
214 92
1 7 6 0 0 4224 0 6 17 0 0 3
484 74
484 147
469 147
1 0 7 0 0 0 0 7 0 0 17 2
389 74
389 147
1 0 8 0 0 0 0 8 0 0 18 2
300 76
300 146
5 0 9 0 0 4096 0 5 0 0 16 2
184 193
184 227
5 0 9 0 0 0 0 13 0 0 16 2
268 194
268 227
5 0 9 0 0 0 0 15 0 0 16 2
357 195
357 227
3 5 9 0 0 4224 0 11 17 0 0 3
160 227
445 227
445 195
3 7 7 0 0 0 0 17 15 0 0 4
415 156
395 156
395 147
381 147
3 7 8 0 0 0 0 15 13 0 0 4
327 156
306 156
306 146
292 146
7 1 2 0 0 0 0 5 9 0 0 3
208 145
214 145
214 76
1 0 10 0 0 4096 0 17 0 0 22 2
445 120
411 120
2 0 10 0 0 0 0 17 0 0 22 2
421 147
411 147
1 4 10 0 0 4224 0 16 17 0 0 3
411 117
411 165
421 165
1 0 11 0 0 4096 0 15 0 0 25 2
357 120
323 120
2 0 11 0 0 0 0 15 0 0 25 2
333 147
323 147
1 4 11 0 0 4224 0 14 15 0 0 3
323 117
323 165
333 165
1 0 12 0 0 4096 0 13 0 0 28 2
268 119
234 119
2 0 12 0 0 0 0 13 0 0 28 2
244 146
234 146
1 4 12 0 0 4224 0 12 13 0 0 3
234 116
234 164
244 164
1 0 13 0 0 4096 0 5 0 0 31 2
184 118
150 118
2 0 13 0 0 0 0 5 0 0 31 2
160 145
150 145
1 4 13 0 0 4224 0 10 5 0 0 3
150 115
150 163
160 163
3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
44 176 72 196
48 180 69 194
3 ___
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 3
42 106 70 126
46 110 67 124
3 ___
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 68
170 275 442 319
174 279 438 311
68 A logic gate implementation of a 
74293 wired as a MOD-16 counter.
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0159882 0 0 0 0.016 0.016
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
