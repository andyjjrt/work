CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 432
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 432
8388626 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 133 194 0 1 11
0 5
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
1 C
-24 -3 -17 5
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 133 138 0 1 11
0 2
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
1 B
-23 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 133 120 0 1 11
0 4
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
1 A
-24 -4 -17 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
8 2-In OR~
219 268 185 0 3 22
0 3 5 6
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
6153 0 0
0
0
8 2-In OR~
219 267 129 0 3 22
0 4 2 7
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
5394 0 0
0
0
9 2-In AND~
219 369 176 0 3 22
0 7 6 8
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7734 0 0
0
0
5 4049~
219 216 176 0 2 22
0 2 3
0
0 0 112 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
15

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0
65 0 0 0 6 2 2 0
1 U
9914 0 0
0
0
14 Logic Display~
6 448 149 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3747 0 0
0
0
8
2 0 2 0 0 4224 0 5 0 0 2 2
254 138
186 138
1 1 2 0 0 0 0 7 2 0 0 4
201 176
186 176
186 138
145 138
2 1 3 0 0 4224 0 7 4 0 0 2
237 176
255 176
1 1 4 0 0 4224 0 5 3 0 0 2
254 120
145 120
2 1 5 0 0 4224 0 4 1 0 0 2
255 194
145 194
2 3 6 0 0 4224 0 6 4 0 0 2
345 185
301 185
1 3 7 0 0 8320 0 6 5 0 0 4
345 167
330 167
330 129
300 129
3 1 8 0 0 4224 0 6 8 0 0 3
390 176
448 176
448 167
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
170 249 186 273
174 253 182 269
1 _
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
468 174 484 198
472 178 480 194
1 _
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
404 188 508 212
408 192 504 208
12 y=(A+B)(B+C)
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 113
58 263 522 307
62 267 518 299
113 Terms A+B and B+C are inputs to an AND gate, and each of 
these two terms is generated from a separate OR gate.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
296 108 320 132
300 112 316 128
2 AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
296 165 320 189
300 169 316 185
2 BC
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
242 158 258 182
246 162 254 178
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
242 150 258 174
246 154 254 170
1 -
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
296 157 312 181
300 161 308 177
1 -
0
2049 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-005 2e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.01 0 0.01 0 0.01 0.01
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 4.81264e-315 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
