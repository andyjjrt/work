CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 8 100 9
4 70 635 430
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 430 635 507
25165842 0
0
6 Title:
5 Name:
0
0
0
16
13 Logic Switch~
5 104 248 0 1 11
0 12
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
2 S1
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 104 232 0 1 11
0 11
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
2 S0
-29 -4 -15 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 486 95 0 1 2
10 5
0
0 0 49264 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
5 SCOPE
12 463 101 0 1 11
0 5
0
0 0 57584 0
1 Z
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
9 3-In AND~
219 333 47 0 4 22
0 9 10 14 18
0
0 0 112 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 1 0
1 U
5394 0 0
0
0
9 3-In AND~
219 333 98 0 4 22
0 8 10 11 17
0
0 0 112 0
6 74LS11
-21 -28 21 -20
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 1 0
1 U
7734 0 0
0
0
9 3-In AND~
219 334 149 0 4 22
0 7 12 13 16
0
0 0 112 0
6 74LS11
-21 -28 21 -20
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 1 0
1 U
9914 0 0
0
0
9 3-In AND~
219 335 200 0 4 22
0 6 12 11 15
0
0 0 112 0
6 74LS11
-21 -28 21 -20
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
3747 0 0
0
0
8 4-In OR~
219 405 123 0 5 22
0 18 17 16 15 5
0
0 0 112 0
4 4072
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0
65 0 0 0 2 1 3 0
1 U
3549 0 0
0
0
9 Inverter~
13 272 70 0 2 22
0 11 14
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
7931 0 0
0
0
9 Inverter~
13 273 168 0 2 22
0 11 13
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
9325 0 0
0
0
9 Inverter~
13 222 117 0 2 22
0 12 10
0
0 0 112 90
6 74LS04
-21 -19 21 -11
3 U4C
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
8903 0 0
0
0
7 Pulser~
4 111 47 0 10 12
0 20 21 9 22 0 0 40 40 39
7
0
0 0 1072 0
0
2 V3
-7 -28 7 -20
4 1kHz
-14 -15 14 -7
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3834 0 0
0
0
7 Pulser~
4 111 98 0 10 12
0 23 24 8 25 0 0 20 20 19
7
0
0 0 1072 0
0
2 V4
-7 -28 7 -20
4 2kHz
-14 -15 14 -7
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3363 0 0
0
0
7 Pulser~
4 111 149 0 10 12
0 26 27 7 28 0 0 15 15 9
8
0
0 0 1072 0
0
2 V5
-7 -28 7 -20
4 3kHz
-14 -15 14 -7
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7668 0 0
0
0
7 Pulser~
4 111 200 0 10 12
0 29 30 6 31 0 0 10 10 9
7
0
0 0 1072 0
0
2 V6
-7 -28 7 -20
4 4kHz
-14 -15 14 -7
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4718 0 0
0
0
26
0 0 1 0 0 4256 0 0 0 0 0 2
517 155
517 234
0 0 2 0 0 4224 0 0 0 0 0 2
468 234
569 234
0 0 3 0 0 4224 0 0 0 0 0 2
469 155
570 155
0 0 4 0 0 4224 0 0 0 0 0 2
469 171
570 171
1 0 5 0 0 4096 0 3 0 0 6 2
486 113
463 113
1 5 5 0 0 8320 0 4 9 0 0 3
463 113
463 123
438 123
1 3 6 0 0 4224 0 8 16 0 0 2
311 191
135 191
1 3 7 0 0 4224 0 7 15 0 0 2
310 140
135 140
1 3 8 0 0 4224 0 6 14 0 0 2
309 89
135 89
1 3 9 0 0 4224 0 5 13 0 0 2
309 38
135 38
2 0 10 0 0 4224 0 6 0 0 19 2
309 98
225 98
3 0 11 0 0 4096 0 6 0 0 17 2
309 107
245 107
2 0 12 0 0 4096 0 7 0 0 18 2
310 149
225 149
3 0 11 0 0 4096 0 8 0 0 17 2
311 209
245 209
2 0 12 0 0 4096 0 8 0 0 18 2
311 200
225 200
1 0 11 0 0 0 0 11 0 0 17 2
258 168
245 168
1 1 11 0 0 8320 0 10 2 0 0 4
257 70
245 70
245 232
116 232
1 1 12 0 0 4224 0 12 1 0 0 3
225 135
225 248
116 248
2 2 10 0 0 0 0 5 12 0 0 3
309 47
225 47
225 99
3 2 13 0 0 8320 0 7 11 0 0 4
310 158
302 158
302 168
294 168
3 2 14 0 0 8320 0 5 10 0 0 4
309 56
301 56
301 70
293 70
4 4 15 0 0 8320 0 8 9 0 0 4
356 200
380 200
380 137
388 137
3 4 16 0 0 4224 0 9 7 0 0 4
388 128
362 128
362 149
355 149
2 4 17 0 0 4224 0 9 6 0 0 4
388 119
362 119
362 98
354 98
4 1 18 0 0 8320 0 5 9 0 0 4
354 47
380 47
380 110
388 110
0 0 19 0 0 4224 0 0 0 0 0 5
299 266
570 266
570 299
299 299
299 266
7
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 23
46 278 238 302
50 282 234 298
23 Four-input multiplexer.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
301 263 567 300
305 267 564 295
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
157 19 181 43
161 23 177 39
2 I0
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
157 70 181 94
161 74 177 90
2 I1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
157 121 181 145
161 125 177 141
2 I2
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
156 172 180 196
160 176 176 192
2 I3
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
469 151 573 255
473 155 569 235
64 S1 S0 Output
0  0   Z=I0
0  1   Z=I1
1  0   Z=I2
1  1   Z=I3
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
267780172 8525888 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 1e-006 2
2
221 112
0 7 0 0 2	0 27 0 0
367 106
0 2 0 0 1	0 27 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 27 0 0
200 112
0 7 0 0 2	0 27 0 0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
