CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 471
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 471
8388626 0
0
6 Title:
5 Name:
0
0
0
46
13 Logic Switch~
5 104 116 0 1 11
0 3
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
2 A3
-30 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 104 133 0 1 11
0 6
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
8 (MSB) A4
-72 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 105 81 0 1 11
0 7
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
2 A2
-30 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 105 63 0 1 11
0 8
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
2 A1
-30 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 105 45 0 1 11
0 9
0
0 0 21616 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
2 A0
-30 -4 -16 4
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5394 0 0
0
0
9 Inverter~
13 432 116 0 2 22
0 3 4
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
7734 0 0
0
0
2 +V
167 164 158 0 1 3
0 5
0
0 0 53616 0
3 +5V
1 -12 22 -4
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9914 0 0
0
0
7 Ground~
168 229 160 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 330 159 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3549 0 0
0
0
7 Ground~
168 430 160 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7931 0 0
0
0
7 74LS138
19 186 206 0 14 29
0 7 8 9 5 6 3 13 12 11
10 14 15 16 17
0
0 0 5232 270
7 74LS138
-25 -61 24 -53
2 U1
-7 -71 7 -63
8 74ALS138
-27 -7 29 1
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
9325 0 0
0
0
7 74LS138
19 286 206 0 14 29
0 7 8 9 3 6 2 37 36 35
34 38 39 40 41
0
0 0 5232 270
7 74LS138
-25 -61 24 -53
2 U2
-7 -71 7 -63
8 74ALS138
-28 -7 28 1
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
8903 0 0
0
0
7 74LS138
19 386 206 0 14 29
0 7 8 9 6 3 2 29 28 27
26 30 31 32 33
0
0 0 5232 270
7 74LS138
-25 -61 24 -53
2 U3
-7 -71 7 -63
8 74ALS138
-27 -7 29 1
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3834 0 0
0
0
7 74LS138
19 486 206 0 14 29
0 7 8 9 6 4 2 21 20 19
18 22 23 24 25
0
0 0 5232 270
7 74LS138
-25 -61 24 -53
2 U4
-7 -71 7 -63
8 74ALS138
-26 -7 30 1
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
14 Logic Display~
6 282 255 0 1 2
10 34
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L9
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7668 0 0
0
0
14 Logic Display~
6 291 255 0 1 2
10 35
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L10
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 300 255 0 1 2
10 36
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L11
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 309 255 0 1 2
10 37
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L12
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6671 0 0
0
0
14 Logic Display~
6 273 255 0 1 2
10 38
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L13
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3789 0 0
0
0
14 Logic Display~
6 264 255 0 1 2
10 39
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L14
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 255 255 0 1 2
10 40
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L15
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3750 0 0
0
0
14 Logic Display~
6 246 255 0 1 2
10 41
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L16
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8778 0 0
0
0
14 Logic Display~
6 382 255 0 1 2
10 26
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L17
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
538 0 0
0
0
14 Logic Display~
6 391 255 0 1 2
10 27
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L18
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6843 0 0
0
0
14 Logic Display~
6 400 255 0 1 2
10 28
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L19
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3136 0 0
0
0
14 Logic Display~
6 409 255 0 1 2
10 29
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L20
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5950 0 0
0
0
14 Logic Display~
6 373 255 0 1 2
10 30
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L21
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5670 0 0
0
0
14 Logic Display~
6 364 255 0 1 2
10 31
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L22
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6828 0 0
0
0
14 Logic Display~
6 355 255 0 1 2
10 32
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L23
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6735 0 0
0
0
14 Logic Display~
6 346 255 0 1 2
10 33
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L24
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8365 0 0
0
0
14 Logic Display~
6 482 255 0 1 2
10 18
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L25
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4132 0 0
0
0
14 Logic Display~
6 491 255 0 1 2
10 19
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L26
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4551 0 0
0
0
14 Logic Display~
6 500 255 0 1 2
10 20
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L27
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3635 0 0
0
0
14 Logic Display~
6 509 255 0 1 2
10 21
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L28
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3973 0 0
0
0
14 Logic Display~
6 473 255 0 1 2
10 22
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L29
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3851 0 0
0
0
14 Logic Display~
6 464 255 0 1 2
10 23
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L30
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8383 0 0
0
0
14 Logic Display~
6 455 255 0 1 2
10 24
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L31
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9334 0 0
0
0
14 Logic Display~
6 446 255 0 1 2
10 25
0
0 0 53360 180
6 100MEG
3 -16 45 -8
3 L32
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7471 0 0
0
0
14 Logic Display~
6 182 255 0 1 2
10 10
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L8
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3334 0 0
0
0
14 Logic Display~
6 191 255 0 1 2
10 11
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L7
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3559 0 0
0
0
14 Logic Display~
6 200 255 0 1 2
10 12
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L6
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
984 0 0
0
0
14 Logic Display~
6 209 255 0 1 2
10 13
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L5
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7557 0 0
0
0
14 Logic Display~
6 173 255 0 1 2
10 14
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L4
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3146 0 0
0
0
14 Logic Display~
6 164 255 0 1 2
10 15
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L3
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5687 0 0
0
0
14 Logic Display~
6 155 255 0 1 2
10 16
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L2
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7939 0 0
0
0
14 Logic Display~
6 146 255 0 1 2
10 17
0
0 0 53360 180
6 100MEG
3 -16 45 -8
2 L1
12 0 26 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3308 0 0
0
0
57
6 0 3 0 0 4112 0 11 0 0 5 2
146 166
146 116
4 0 3 0 0 4112 0 12 0 0 5 2
264 172
264 116
5 0 3 0 0 16 0 13 0 0 5 2
355 166
355 116
2 5 4 0 0 8336 0 6 14 0 0 3
453 116
455 116
455 166
1 1 3 0 0 4240 0 1 6 0 0 2
116 116
417 116
1 4 5 0 0 4240 0 7 11 0 0 2
164 167
164 172
1 6 2 0 0 4240 0 8 12 0 0 3
229 154
246 154
246 166
1 6 2 0 0 16 0 9 13 0 0 3
330 153
346 153
346 166
1 6 2 0 0 16 0 10 14 0 0 3
430 154
446 154
446 166
5 0 6 0 0 4112 0 11 0 0 13 2
155 166
155 133
5 0 6 0 0 16 0 12 0 0 13 2
255 166
255 133
4 0 6 0 0 4112 0 13 0 0 13 2
364 172
364 133
1 4 6 0 0 4240 0 2 14 0 0 3
116 133
464 133
464 172
1 0 7 0 0 4112 0 11 0 0 17 2
209 172
209 81
1 0 7 0 0 16 0 12 0 0 17 2
309 172
309 81
1 0 7 0 0 16 0 13 0 0 17 2
409 172
409 81
1 1 7 0 0 4240 0 3 14 0 0 3
117 81
509 81
509 172
2 0 8 0 0 4112 0 11 0 0 21 2
200 172
200 63
2 0 8 0 0 16 0 12 0 0 21 2
300 172
300 63
2 0 8 0 0 16 0 13 0 0 21 2
400 172
400 63
1 2 8 0 0 4240 0 4 14 0 0 3
117 63
500 63
500 172
3 0 9 0 0 4112 0 11 0 0 25 2
191 172
191 45
3 0 9 0 0 16 0 12 0 0 25 2
291 172
291 45
3 0 9 0 0 16 0 13 0 0 25 2
391 172
391 45
1 3 9 0 0 4240 0 5 14 0 0 3
117 45
491 45
491 172
1 10 10 0 0 4240 0 39 11 0 0 2
182 241
182 242
1 9 11 0 0 4240 0 40 11 0 0 2
191 241
191 242
1 8 12 0 0 4240 0 41 11 0 0 2
200 241
200 242
1 7 13 0 0 4240 0 42 11 0 0 2
209 241
209 242
1 11 14 0 0 4240 0 43 11 0 0 2
173 241
173 242
1 12 15 0 0 4240 0 44 11 0 0 2
164 241
164 242
1 13 16 0 0 4240 0 45 11 0 0 2
155 241
155 242
1 14 17 0 0 4240 0 46 11 0 0 2
146 241
146 242
1 10 18 0 0 4240 0 31 14 0 0 2
482 241
482 242
1 9 19 0 0 4240 0 32 14 0 0 2
491 241
491 242
1 8 20 0 0 4240 0 33 14 0 0 2
500 241
500 242
1 7 21 0 0 4240 0 34 14 0 0 2
509 241
509 242
1 11 22 0 0 4240 0 35 14 0 0 2
473 241
473 242
1 12 23 0 0 4240 0 36 14 0 0 2
464 241
464 242
1 13 24 0 0 4240 0 37 14 0 0 2
455 241
455 242
1 14 25 0 0 4240 0 38 14 0 0 2
446 241
446 242
1 10 26 0 0 4240 0 23 13 0 0 2
382 241
382 242
1 9 27 0 0 4240 0 24 13 0 0 2
391 241
391 242
1 8 28 0 0 4240 0 25 13 0 0 2
400 241
400 242
1 7 29 0 0 4240 0 26 13 0 0 2
409 241
409 242
1 11 30 0 0 4240 0 27 13 0 0 2
373 241
373 242
1 12 31 0 0 4240 0 28 13 0 0 2
364 241
364 242
1 13 32 0 0 4240 0 29 13 0 0 2
355 241
355 242
1 14 33 0 0 4240 0 30 13 0 0 2
346 241
346 242
1 10 34 0 0 4240 0 15 12 0 0 2
282 241
282 242
1 9 35 0 0 4240 0 16 12 0 0 2
291 241
291 242
1 8 36 0 0 4240 0 17 12 0 0 2
300 241
300 242
1 7 37 0 0 4240 0 18 12 0 0 2
309 241
309 242
1 11 38 0 0 4240 0 19 12 0 0 2
273 241
273 242
1 12 39 0 0 4240 0 20 12 0 0 2
264 241
264 242
1 13 40 0 0 4240 0 21 12 0 0 2
255 241
255 242
1 14 41 0 0 4240 0 22 12 0 0 2
246 241
246 242
13
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
135 271 219 291
139 275 216 289
11 O0-------O7
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
336 271 420 291
340 275 417 289
11 O16-----O23
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
235 271 319 291
239 275 316 289
11 O8------O15
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 11
436 271 520 291
440 275 517 289
11 O24-----O31
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
135 259 149 279
139 263 146 277
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
198 259 212 279
202 263 209 277
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
235 259 249 279
239 263 246 277
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
291 259 305 279
295 263 302 277
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
336 259 350 279
340 263 347 277
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
392 259 406 279
396 263 403 277
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
436 259 450 279
440 263 447 277
1 _
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
492 259 506 279
496 263 503 277
1 _
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 41
144 323 480 347
148 327 476 343
41 Four 74ALS138s forming a 1-of-32 decoder.
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
267780172 8525888 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
9.98039 0 5.4 0 10 10
12401 0
4 1e-006 2
2
221 112
0 7 0 0 2	0 58 0 0
367 106
0 2 0 0 1	0 58 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
9.98039 0 5.4 0 10 10
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 58 0 0
200 112
0 7 0 0 2	0 58 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
