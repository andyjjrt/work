CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 375
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 375 635 485
25165842 0
0
6 Title:
5 Name:
0
0
0
5
5 SCOPE
12 244 82 0 1 11
0 5
0
0 0 57584 0
1 A
-4 -4 3 4
2 U2
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
5 SCOPE
12 284 82 0 1 11
0 4
0
0 0 57584 0
1 B
-4 -4 3 4
2 U3
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 391 83 0 1 11
0 3
0
0 0 57584 0
1 x
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
9 Data Seq~
170 179 82 0 17 18
0 6 7 8 9 10 11 4 5 12
13 18 1 20 10 5 0 33
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
6153 0 0
0
0
AAAAABACADACADACADAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAABAAAB
9 2-In AND~
219 333 127 0 3 22
0 5 4 3
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5394 0 0
0
0
6
0 0 2 0 0 4224 0 0 0 0 0 5
305 206
574 206
574 239
305 239
305 206
1 3 3 0 0 8320 0 3 5 0 0 3
391 95
391 127
354 127
1 0 4 0 0 4096 0 2 0 0 5 2
284 94
284 109
1 0 5 0 0 4096 0 1 0 0 6 2
244 94
244 118
7 2 4 0 0 4224 0 4 5 0 0 4
211 109
284 109
284 136
309 136
8 1 5 0 0 4224 0 4 5 0 0 2
211 118
309 118
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
71 212 215 236
75 216 211 232
17 2-input AND gate.
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
307 203 573 240
311 207 570 235
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 2
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 2e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.0022 0.0008 30 -30 0.003 0.003
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
