CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
4 70 635 458
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
4 70 635 458
8912914 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 67 141 0 1 11
0 8
0
0 0 21616 0
2 0V
-6 -16 8 -8
4 VIN1
-39 -4 -11 4
1 B
-22 -5 -15 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 66 82 0 1 11
0 9
0
0 0 21616 0
2 0V
-6 -16 8 -8
3 VIN
-36 -4 -15 4
1 A
-23 -5 -16 3
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
7 Ground~
168 364 178 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
11 Multimeter~
205 339 144 0 21 21
0 7 12 13 2 0 0 0 0 0
78 79 32 68 65 84 65 32 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM1
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
6153 0 0
0
0
12 N-EMOS 3T:A~
219 266 213 0 3 7
0 7 8 2
0
0 0 1104 512
4 NMOS
18 0 46 8
2 Q2
18 -5 32 3
2 Q2
-36 -5 -22 3
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 1 2 3 1 2 3 0
77 0 0 0 0 0 0 0
1 Q
5394 0 0
0
0
12 N-EMOS 3T:A~
219 182 213 0 3 7
0 7 9 2
0
0 0 1104 0
4 NMOS
18 0 46 8
2 Q6
18 -5 32 3
2 Q2
18 -5 32 3
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 1 2 3 1 2 3 0
77 0 0 0 0 0 0 0
1 Q
7734 0 0
0
0
2 +V
167 221 43 0 1 3
0 11
0
0 0 54384 0
2 5V
-7 -22 7 -14
2 V3
-7 -32 7 -24
4 +VDD
-12 -14 16 -6
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9914 0 0
0
0
7 Ground~
168 221 257 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3747 0 0
0
0
12 P-EMOS 3T:A~
219 215 91 0 3 7
0 10 9 11
0
0 0 1104 692
4 PMOS
18 0 46 8
2 Q5
18 -5 32 3
2 Q1
18 -5 32 3
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 2 3 1 2 3 1 0
109 0 0 0 0 0 0 0
1 Q
3549 0 0
0
0
12 P-EMOS 3T:A~
219 215 150 0 3 7
0 7 8 10
0
0 0 1104 692
4 PMOS
18 0 46 8
2 Q1
18 -5 32 3
2 Q1
18 -5 32 3
0
17 %D %1 %2 %3 %3 %M
0
0
0
7

0 2 3 1 2 3 1 0
109 0 0 0 0 0 0 0
1 Q
7931 0 0
0
0
17
0 0 1 0 0 4272 0 0 0 4 3 2
505 141
505 220
0 0 3 0 0 4240 0 0 0 0 0 2
461 145
461 216
0 0 4 0 0 4240 0 0 0 0 0 2
424 220
547 220
0 0 5 0 0 4240 0 0 0 0 0 2
423 141
546 141
0 0 6 0 0 4240 0 0 0 0 0 2
423 156
546 156
0 1 7 0 0 4224 0 0 4 11 0 3
221 175
314 175
314 167
2 0 8 0 0 12416 0 5 0 0 9 5
280 222
289 222
289 275
110 275
110 141
2 0 9 0 0 8320 0 6 0 0 10 3
164 222
137 222
137 82
1 2 8 0 0 0 0 1 10 0 0 2
79 141
197 141
1 2 9 0 0 0 0 2 9 0 0 2
78 82
197 82
1 0 7 0 0 0 0 10 0 0 14 2
221 168
221 187
1 0 2 0 0 4096 0 8 0 0 13 2
221 251
221 239
3 3 2 0 0 8320 0 6 5 0 0 4
188 231
188 239
256 239
256 231
1 1 7 0 0 0 0 6 5 0 0 4
188 195
188 187
256 187
256 195
1 3 10 0 0 4224 0 9 10 0 0 2
221 109
221 132
1 3 11 0 0 4224 0 7 9 0 0 2
221 52
221 73
1 4 2 0 0 0 0 3 4 0 0 2
364 172
364 167
4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
239 310 359 334
243 314 355 330
14 CMOS NOR gate.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
265 141 297 165
269 145 293 161
3 ___
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
249 156 297 180
253 160 293 176
5 X=A+B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 78
421 137 557 241
425 141 553 221
78  A    B     X
LOW  LOW   HIGH
LOW  HIGH  LOW
HIGH LOW   LOW
HIGH HIGH  LOW
0
1 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
-1235812058 1210432 100 100 0 0
77 66 587 246
420 103 581 173
587 66
77 66
587 66
587 246
0 0
0.003 0 5.4 0 0.003 5.4
12401 0
4 2 2
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
