CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 5 100 9
4 70 635 430
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 430 635 709
25165842 0
0
6 Title:
5 Name:
0
0
0
34
9 Inverter~
13 360 159 0 2 22
0 12 15
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U4C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
8953 0 0
0
0
9 Inverter~
13 359 117 0 2 22
0 2 13
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U4B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
4441 0 0
0
0
9 Inverter~
13 358 62 0 2 22
0 11 14
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
3618 0 0
0
0
9 3-In AND~
219 467 282 0 4 22
0 11 2 12 3
0
0 0 1120 0
6 74LS11
-21 -28 21 -20
3 U3B
-12 -25 9 -17
1 7
-6 -4 1 4
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 3 0
1 U
6153 0 0
0
0
9 3-In AND~
219 467 249 0 4 22
0 14 2 12 4
0
0 0 1120 0
6 74LS11
-21 -28 21 -20
3 U3A
-12 -25 9 -17
1 6
-6 -4 1 4
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 3 0
1 U
5394 0 0
0
0
9 3-In AND~
219 467 216 0 4 22
0 11 13 12 5
0
0 0 1120 0
6 74LS11
-21 -28 21 -20
3 U2C
-12 -25 9 -17
1 5
-6 -4 1 4
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 2 0
1 U
7734 0 0
0
0
9 3-In AND~
219 467 183 0 4 22
0 14 13 12 6
0
0 0 1120 0
6 74LS11
-21 -28 21 -20
3 U2B
-12 -25 9 -17
1 4
-6 -4 1 4
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 2 0
1 U
9914 0 0
0
0
9 3-In AND~
219 467 150 0 4 22
0 11 2 15 7
0
0 0 1120 0
6 74LS11
-21 -28 21 -20
3 U2A
-12 -25 9 -17
1 3
-6 -4 1 4
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
3747 0 0
0
0
9 3-In AND~
219 467 117 0 4 22
0 14 2 15 8
0
0 0 1120 0
6 74LS11
-21 -28 21 -20
3 U1C
-12 -25 9 -17
1 2
-6 -4 1 4
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 1 0
1 U
3549 0 0
0
0
9 3-In AND~
219 467 84 0 4 22
0 11 13 15 9
0
0 0 1120 0
6 74LS11
-21 -28 21 -20
3 U1B
-12 -25 9 -17
1 1
-6 -4 1 4
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 1 0
1 U
7931 0 0
0
0
9 3-In AND~
219 467 51 0 4 22
0 14 13 15 10
0
0 0 1120 0
6 74LS11
-21 -28 21 -20
3 U1A
-12 -25 9 -17
1 0
-6 -4 1 4
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 1 0
1 U
9325 0 0
0
0
9 Data Seq~
170 121 107 0 17 18
0 17 18 19 20 21 12 2 11 22
23 1 1 8 5 6 0 33
0
0 0 4192 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
8903 0 0
0
0
AAAAABACADAEAFAGAHAAABACADAEAFAGAHAAABACADAEAFAGAHAAABACADAEAFAGAH
5 SCOPE
12 279 87 0 1 11
0 11
0
0 0 57568 0
1 A
-4 -4 3 4
2 U7
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3834 0 0
0
0
5 SCOPE
12 229 87 0 1 11
0 2
0
0 0 57568 0
1 B
-4 -4 3 4
2 U6
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3363 0 0
0
0
5 SCOPE
12 179 87 0 1 11
0 12
0
0 0 57568 0
1 C
-4 -4 3 4
2 U5
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
7668 0 0
0
0
14 Logic Display~
6 202 81 0 1 2
10 12
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4718 0 0
0
0
14 Logic Display~
6 252 81 0 1 2
10 2
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3874 0 0
0
0
14 Logic Display~
6 302 81 0 1 2
10 11
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6671 0 0
0
0
5 SCOPE
12 502 38 0 1 11
0 10
0
0 0 57568 0
2 O0
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3789 0 0
0
0
14 Logic Display~
6 526 32 0 1 2
10 10
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 526 65 0 1 2
10 9
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3750 0 0
0
0
5 SCOPE
12 502 71 0 1 11
0 9
0
0 0 57568 0
2 O1
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8778 0 0
0
0
14 Logic Display~
6 526 98 0 1 2
10 8
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
538 0 0
0
0
5 SCOPE
12 502 104 0 1 11
0 8
0
0 0 57568 0
2 O2
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6843 0 0
0
0
14 Logic Display~
6 526 131 0 1 2
10 7
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3136 0 0
0
0
5 SCOPE
12 502 137 0 1 11
0 7
0
0 0 57568 0
2 O3
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
5950 0 0
0
0
14 Logic Display~
6 526 164 0 1 2
10 6
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
5 SCOPE
12 502 170 0 1 11
0 6
0
0 0 57568 0
2 O4
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6828 0 0
0
0
14 Logic Display~
6 526 197 0 1 2
10 5
0
0 0 53360 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
5 SCOPE
12 502 203 0 1 11
0 5
0
0 0 57568 0
2 O5
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
8365 0 0
0
0
14 Logic Display~
6 526 230 0 1 2
10 4
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4132 0 0
0
0
5 SCOPE
12 502 236 0 1 11
0 4
0
0 0 57568 0
2 O6
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4551 0 0
0
0
14 Logic Display~
6 526 263 0 1 2
10 3
0
0 0 53360 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3635 0 0
0
0
5 SCOPE
12 502 269 0 1 11
0 3
0
0 0 57568 0
2 O7
-8 -4 6 4
2 U8
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3973 0 0
0
0
50
0 0 16 0 0 16 0 0 0 0 0 5
17 244
288 244
288 275
17 275
17 244
0 7 2 0 0 4224 0 0 12 48 0 2
425 134
153 134
1 0 3 0 0 8320 0 33 0 0 4 3
526 281
526 282
502 282
1 4 3 0 0 0 0 34 4 0 0 3
502 281
502 282
488 282
1 0 4 0 0 8320 0 31 0 0 6 3
526 248
526 249
502 249
1 4 4 0 0 0 0 32 5 0 0 3
502 248
502 249
488 249
1 0 5 0 0 8320 0 29 0 0 8 3
526 215
526 216
502 216
1 4 5 0 0 0 0 30 6 0 0 3
502 215
502 216
488 216
1 0 6 0 0 8320 0 27 0 0 10 3
526 182
526 183
502 183
1 4 6 0 0 0 0 28 7 0 0 3
502 182
502 183
488 183
1 0 7 0 0 8320 0 25 0 0 12 3
526 149
526 150
502 150
1 4 7 0 0 0 0 26 8 0 0 3
502 149
502 150
488 150
1 0 8 0 0 8320 0 23 0 0 14 3
526 116
526 117
502 117
1 4 8 0 0 0 0 24 9 0 0 3
502 116
502 117
488 117
1 0 9 0 0 8320 0 21 0 0 16 3
526 83
526 84
502 84
1 4 9 0 0 0 0 22 10 0 0 3
502 83
502 84
488 84
1 0 10 0 0 8320 0 20 0 0 18 3
526 50
526 51
502 51
1 4 10 0 0 0 0 19 11 0 0 3
502 50
502 51
488 51
1 0 11 0 0 4096 0 18 0 0 29 2
302 99
302 143
1 0 11 0 0 0 0 13 0 0 29 2
279 99
279 143
1 0 2 0 0 0 0 17 0 0 2 2
252 99
252 134
1 0 2 0 0 0 0 14 0 0 2 2
229 99
229 134
1 0 12 0 0 4096 0 16 0 0 28 2
202 99
202 125
1 0 12 0 0 0 0 15 0 0 28 2
179 99
179 125
1 0 12 0 0 8192 0 1 0 0 28 3
345 159
334 159
334 192
1 0 2 0 0 0 0 2 0 0 2 3
344 117
334 117
334 134
1 0 11 0 0 0 0 3 0 0 29 3
343 62
334 62
334 84
0 6 12 0 0 12416 0 0 12 49 0 4
435 192
313 192
313 125
153 125
0 8 11 0 0 12288 0 0 12 46 0 4
405 84
322 84
322 143
153 143
3 0 12 0 0 0 0 5 0 0 49 2
443 258
435 258
2 0 2 0 0 0 0 5 0 0 48 2
443 249
425 249
3 0 12 0 0 0 0 6 0 0 49 2
443 225
435 225
1 0 11 0 0 0 0 6 0 0 46 2
443 207
405 207
2 0 13 0 0 4096 0 7 0 0 47 2
443 183
415 183
1 0 14 0 0 4096 0 7 0 0 45 2
443 174
395 174
2 0 2 0 0 0 0 8 0 0 48 2
443 150
425 150
1 0 11 0 0 0 0 8 0 0 46 2
443 141
405 141
3 0 15 0 0 4096 0 9 0 0 50 2
443 126
435 126
1 0 14 0 0 0 0 9 0 0 45 2
443 108
395 108
3 0 15 0 0 0 0 10 0 0 50 2
443 93
435 93
2 0 13 0 0 0 0 10 0 0 47 2
443 84
415 84
2 0 14 0 0 0 0 3 0 0 45 2
379 62
395 62
2 0 13 0 0 4096 0 2 0 0 47 2
380 117
415 117
2 0 15 0 0 4096 0 1 0 0 50 2
381 159
435 159
1 1 14 0 0 8320 0 11 5 0 0 4
443 42
395 42
395 240
443 240
1 1 11 0 0 8320 0 10 4 0 0 4
443 75
405 75
405 273
443 273
2 2 13 0 0 8320 0 11 6 0 0 4
443 51
415 51
415 216
443 216
2 2 2 0 0 0 0 9 4 0 0 4
443 117
425 117
425 282
443 282
3 3 12 0 0 0 0 7 4 0 0 4
443 192
435 192
435 291
443 291
3 3 15 0 0 8320 0 11 8 0 0 4
443 60
435 60
435 159
443 159
2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
19 241 285 278
23 245 282 273
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 1
-13 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 37
9 285 313 309
13 289 309 305
37 3-line-to-8-line (or 1-of-8) decoder.
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 10 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
267780172 8525888 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
9.98039 0 5.4 0 10 10
12401 0
4 1e-006 2
2
221 112
0 7 0 0 2	0 51 0 0
367 106
0 2 0 0 1	0 51 0 0
1208353588 8788032 100 100 0 0
77 66 587 216
4 430 635 712
586 66
77 66
587 66
587 216
0 0
0.00214706 0.000547058 4.8 1.70667 0.003 0.003
12401 0
4 1e-006 2
2
331 106
0 2 0 0 1	0 51 0 0
200 112
0 7 0 0 2	0 51 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
