CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
4 70 635 393
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
65 C:\Program Files\MicroCode Engineering\CircuitMaker 6 Pro\BOM.DAT
0 7
3 393 635 502
25165842 0
0
6 Title:
5 Name:
0
0
0
5
5 4011~
219 210 135 0 3 22
0 7 6 8
0
0 0 112 0
4 4011
-7 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 589827
65 0 0 0 4 1 1 0
1 U
8953 0 0
0
0
5 SCOPE
12 132 80 0 1 11
0 7
0
0 0 57584 0
1 A
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
5 SCOPE
12 167 80 0 1 11
0 6
0
0 0 57584 0
1 B
-4 -4 3 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
3618 0 0
0
0
5 SCOPE
12 265 80 0 1 11
0 8
0
0 0 57584 0
3 Out
-11 -4 10 4
2 U4
-8 -14 6 -6
0
0
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
0
6153 0 0
0
0
9 Data Seq~
170 71 90 0 17 18
0 9 10 11 12 13 14 6 7 15
16 1 1 60 10 11 0 65
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -44 10 -36
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
5394 0 0
0
0
AAACACADADACAAABABABABADADACACADADABABAAAAAAAAAAAAAAAAAAAAAAAAAAAAACACACACACACAC
ACACACACACACACACACACACACACACACACACACACACACACACACAC
10
0 0 2 0 0 4224 0 0 0 0 0 5
310 222
579 222
579 255
310 255
310 222
0 0 1 0 0 4256 0 0 0 5 3 2
454 58
454 144
0 0 3 0 0 4224 0 0 0 0 0 2
394 144
486 144
0 0 4 0 0 4224 0 0 0 0 0 2
394 77
486 77
0 0 5 0 0 4224 0 0 0 0 0 2
394 58
486 58
1 0 6 0 0 4096 0 3 0 0 9 2
167 92
167 144
1 0 7 0 0 4096 0 2 0 0 8 2
132 92
132 126
1 8 7 0 0 4224 0 1 5 0 0 2
186 126
103 126
2 7 6 0 0 4224 0 1 5 0 0 4
186 144
118 144
118 117
103 117
3 1 8 0 0 8320 0 1 4 0 0 3
237 135
265 135
265 92
6
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 64
312 219 578 256
316 223 575 251
64 Select 'Simulation > Digital Options'
Set 'X Magnification' = 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
228 146 268 170
232 150 264 166
4 x=AB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
245 131 269 155
249 135 265 151
2 __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
455 44 487 68
459 48 483 64
3  __
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 59
391 58 487 162
395 62 483 142
59 A   B    AB
0   0    1
0   1    1
1   0    1
1   1    0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 26
28 230 244 254
32 234 240 250
26 NAND gate and truth table.
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 6e-005 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
449119056 1210432 100 100 0 0
0 0 0 0
11 95 172 165
0 0
0 0
0 0
0 0
0 0
0.00405882 0.00269412 4.2 1.60756e-314 0.006 0.006
12401 0
4 3 10000
0
65864252 8550464 100 100 0 0
77 66 587 246
4 405 625 740
587 66
77 66
587 66
587 246
0 0
0.005 0 6 -6 0.005 0.005
12401 0
4 0.001 2e+012
0
0 0 100 100 0 0
77 66 587 216
0 0 0 0
587 66
77 66
587 66
587 216
0 0
400 100 400 100 300 300
12385 0
0 100000 200000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
